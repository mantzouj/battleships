
module DE2_Audio_Example (
	// Inputs
	CLOCK_50,
	CLOCK_27,
	KEY,

	AUD_ADCDAT,

	// Bidirectionals
	AUD_BCLK,
	AUD_ADCLRCK,
	AUD_DACLRCK,

	I2C_SDAT,

	// Outputs
	AUD_XCK,
	AUD_DACDAT,

	I2C_SCLK,
	SW,
	test
);

/*****************************************************************************
 *                           Parameter Declarations                          *
 *****************************************************************************/


/*****************************************************************************
 *                             Port Declarations                             *
 *****************************************************************************/
// Inputs
input				CLOCK_50;
input				CLOCK_27;
input		[3:0]	KEY;
input				SW;
input				AUD_ADCDAT;

// Bidirectionals
inout				AUD_BCLK;
inout				AUD_ADCLRCK;
inout				AUD_DACLRCK;

inout				I2C_SDAT;

// Outputs
output				AUD_XCK;
output				AUD_DACDAT;
output				test;

output				I2C_SCLK;

/*****************************************************************************
 *                 Internal Wires and Registers Declarations                 *
 *****************************************************************************/
// Internal Wires
wire				audio_in_available;
wire		[31:0]	left_channel_audio_in;
wire		[31:0]	right_channel_audio_in;
wire				read_audio_in;

wire				audio_out_allowed;
wire		[31:0]	left_channel_audio_out;
wire		[31:0]	right_channel_audio_out;
wire				write_audio_out;

// Internal Registers

reg [16:0] delay_cnt;
reg signed [31:0] sound1;
reg [12:0] counter;
reg snd, start, testi;

// State Machine Registers

/*****************************************************************************
 *                         Finite State Machine(s)                           *
 *****************************************************************************/


/*****************************************************************************
 *                             Sequential Logic                              *
 *****************************************************************************/

always @(posedge CLOCK_50) begin
	if(SW == 0) begin
		counter <= 13'd0;
		delay_cnt <= 17'd0;
		testi <= 1'b1;
	end else start <= 1'b1;
	
	if (start == 1) begin
	
	if(delay_cnt == 8000) begin
		delay_cnt <= 17'd0;
		counter <= counter + 13'd1;
		case (counter)
	0: sound1 <=  0;
	1: sound1 <=  0;
	2: sound1 <=  0;
	3: sound1 <=  0;
	4: sound1 <=  -92;
	5: sound1 <=  92;
	6: sound1 <=  -244;
	7: sound1 <=  336;
	8: sound1 <=  -732;
	9: sound1 <=  1099;
	10: sound1 <=  -2441;
	11: sound1 <=  10895;
	12: sound1 <=  31586;
	13: sound1 <=  27985;
	14: sound1 <=  29602;
	15: sound1 <=  28839;
	16: sound1 <=  29724;
	17: sound1 <=  29297;
	18: sound1 <=  29205;
	19: sound1 <=  29541;
	20: sound1 <=  29633;
	21: sound1 <=  28992;
	22: sound1 <=  29572;
	23: sound1 <=  29327;
	24: sound1 <=  28809;
	25: sound1 <=  28992;
	26: sound1 <=  29419;
	27: sound1 <=  29388;
	28: sound1 <=  29419;
	29: sound1 <=  29358;
	30: sound1 <=  29602;
	31: sound1 <=  29510;
	32: sound1 <=  29449;
	33: sound1 <=  28992;
	34: sound1 <=  29144;
	35: sound1 <=  29510;
	36: sound1 <=  29236;
	37: sound1 <=  28839;
	38: sound1 <=  28809;
	39: sound1 <=  29510;
	40: sound1 <=  29114;
	41: sound1 <=  29022;
	42: sound1 <=  29114;
	43: sound1 <=  29449;
	44: sound1 <=  29694;
	45: sound1 <=  28839;
	46: sound1 <=  28961;
	47: sound1 <=  29022;
	48: sound1 <=  29144;
	49: sound1 <=  28992;
	50: sound1 <=  29083;
	51: sound1 <=  29236;
	52: sound1 <=  29144;
	53: sound1 <=  28748;
	54: sound1 <=  28992;
	55: sound1 <=  29022;
	56: sound1 <=  29236;
	57: sound1 <=  29480;
	58: sound1 <=  29022;
	59: sound1 <=  29053;
	60: sound1 <=  29266;
	61: sound1 <=  29053;
	62: sound1 <=  29449;
	63: sound1 <=  29724;
	64: sound1 <=  29266;
	65: sound1 <=  29297;
	66: sound1 <=  29297;
	67: sound1 <=  29297;
	68: sound1 <=  29114;
	69: sound1 <=  29083;
	70: sound1 <=  29266;
	71: sound1 <=  29236;
	72: sound1 <=  29297;
	73: sound1 <=  29419;
	74: sound1 <=  28748;
	75: sound1 <=  29205;
	76: sound1 <=  29266;
	77: sound1 <=  29358;
	78: sound1 <=  28992;
	79: sound1 <=  29114;
	80: sound1 <=  29358;
	81: sound1 <=  29114;
	82: sound1 <=  29205;
	83: sound1 <=  29205;
	84: sound1 <=  29510;
	85: sound1 <=  29388;
	86: sound1 <=  29266;
	87: sound1 <=  28961;
	88: sound1 <=  28839;
	89: sound1 <=  29053;
	90: sound1 <=  29114;
	91: sound1 <=  28656;
	92: sound1 <=  29175;
	93: sound1 <=  29022;
	94: sound1 <=  28900;
	95: sound1 <=  28992;
	96: sound1 <=  29022;
	97: sound1 <=  28900;
	98: sound1 <=  29144;
	99: sound1 <=  29144;
	100: sound1 <=  28961;
	101: sound1 <=  29053;
	102: sound1 <=  29358;
	103: sound1 <=  29449;
	104: sound1 <=  29144;
	105: sound1 <=  28992;
	106: sound1 <=  29083;
	107: sound1 <=  28656;
	108: sound1 <=  29053;
	109: sound1 <=  28961;
	110: sound1 <=  28870;
	111: sound1 <=  29236;
	112: sound1 <=  28809;
	113: sound1 <=  29083;
	114: sound1 <=  29327;
	115: sound1 <=  29327;
	116: sound1 <=  28809;
	117: sound1 <=  29266;
	118: sound1 <=  29510;
	119: sound1 <=  29083;
	120: sound1 <=  29175;
	121: sound1 <=  29633;
	122: sound1 <=  29572;
	123: sound1 <=  29083;
	124: sound1 <=  28900;
	125: sound1 <=  29114;
	126: sound1 <=  29083;
	127: sound1 <=  29541;
	128: sound1 <=  29327;
	129: sound1 <=  29266;
	130: sound1 <=  29572;
	131: sound1 <=  29785;
	132: sound1 <=  29846;
	133: sound1 <=  29663;
	134: sound1 <=  29297;
	135: sound1 <=  29541;
	136: sound1 <=  29449;
	137: sound1 <=  29236;
	138: sound1 <=  29419;
	139: sound1 <=  29297;
	140: sound1 <=  29144;
	141: sound1 <=  29266;
	142: sound1 <=  29236;
	143: sound1 <=  29205;
	144: sound1 <=  29175;
	145: sound1 <=  29083;
	146: sound1 <=  28931;
	147: sound1 <=  28931;
	148: sound1 <=  29144;
	149: sound1 <=  29297;
	150: sound1 <=  29022;
	151: sound1 <=  29297;
	152: sound1 <=  29053;
	153: sound1 <=  29053;
	154: sound1 <=  29419;
	155: sound1 <=  29755;
	156: sound1 <=  29266;
	157: sound1 <=  29327;
	158: sound1 <=  29236;
	159: sound1 <=  28992;
	160: sound1 <=  29266;
	161: sound1 <=  29205;
	162: sound1 <=  29205;
	163: sound1 <=  29053;
	164: sound1 <=  29266;
	165: sound1 <=  29175;
	166: sound1 <=  29144;
	167: sound1 <=  29297;
	168: sound1 <=  29083;
	169: sound1 <=  29358;
	170: sound1 <=  29419;
	171: sound1 <=  29694;
	172: sound1 <=  29663;
	173: sound1 <=  29236;
	174: sound1 <=  29663;
	175: sound1 <=  29572;
	176: sound1 <=  29297;
	177: sound1 <=  29388;
	178: sound1 <=  29633;
	179: sound1 <=  28992;
	180: sound1 <=  29633;
	181: sound1 <=  29694;
	182: sound1 <=  29602;
	183: sound1 <=  29602;
	184: sound1 <=  28992;
	185: sound1 <=  29083;
	186: sound1 <=  29327;
	187: sound1 <=  29419;
	188: sound1 <=  29633;
	189: sound1 <=  29388;
	190: sound1 <=  29083;
	191: sound1 <=  29022;
	192: sound1 <=  29449;
	193: sound1 <=  29449;
	194: sound1 <=  29297;
	195: sound1 <=  29175;
	196: sound1 <=  29205;
	197: sound1 <=  29510;
	198: sound1 <=  29083;
	199: sound1 <=  29266;
	200: sound1 <=  28992;
	201: sound1 <=  28625;
	202: sound1 <=  29022;
	203: sound1 <=  28870;
	204: sound1 <=  28931;
	205: sound1 <=  29022;
	206: sound1 <=  28931;
	207: sound1 <=  29205;
	208: sound1 <=  29022;
	209: sound1 <=  29114;
	210: sound1 <=  29114;
	211: sound1 <=  29358;
	212: sound1 <=  29175;
	213: sound1 <=  29083;
	214: sound1 <=  28717;
	215: sound1 <=  29022;
	216: sound1 <=  29205;
	217: sound1 <=  28778;
	218: sound1 <=  28717;
	219: sound1 <=  28900;
	220: sound1 <=  28931;
	221: sound1 <=  28992;
	222: sound1 <=  29083;
	223: sound1 <=  28992;
	224: sound1 <=  29053;
	225: sound1 <=  29175;
	226: sound1 <=  29114;
	227: sound1 <=  28839;
	228: sound1 <=  29053;
	229: sound1 <=  29358;
	230: sound1 <=  28870;
	231: sound1 <=  28778;
	232: sound1 <=  28931;
	233: sound1 <=  29083;
	234: sound1 <=  28992;
	235: sound1 <=  28992;
	236: sound1 <=  28961;
	237: sound1 <=  28992;
	238: sound1 <=  29144;
	239: sound1 <=  29419;
	240: sound1 <=  29144;
	241: sound1 <=  29236;
	242: sound1 <=  29480;
	243: sound1 <=  28625;
	244: sound1 <=  28778;
	245: sound1 <=  28931;
	246: sound1 <=  29083;
	247: sound1 <=  29053;
	248: sound1 <=  29144;
	249: sound1 <=  28870;
	250: sound1 <=  28931;
	251: sound1 <=  29236;
	252: sound1 <=  29053;
	253: sound1 <=  28870;
	254: sound1 <=  29205;
	255: sound1 <=  29449;
	256: sound1 <=  29114;
	257: sound1 <=  28961;
	258: sound1 <=  29358;
	259: sound1 <=  29053;
	260: sound1 <=  29053;
	261: sound1 <=  29633;
	262: sound1 <=  29266;
	263: sound1 <=  29358;
	264: sound1 <=  29236;
	265: sound1 <=  28931;
	266: sound1 <=  29419;
	267: sound1 <=  29205;
	268: sound1 <=  29236;
	269: sound1 <=  29175;
	270: sound1 <=  29785;
	271: sound1 <=  29602;
	272: sound1 <=  29266;
	273: sound1 <=  29419;
	274: sound1 <=  29755;
	275: sound1 <=  29175;
	276: sound1 <=  29022;
	277: sound1 <=  28992;
	278: sound1 <=  29419;
	279: sound1 <=  29175;
	280: sound1 <=  29114;
	281: sound1 <=  29266;
	282: sound1 <=  28961;
	283: sound1 <=  29297;
	284: sound1 <=  29602;
	285: sound1 <=  29297;
	286: sound1 <=  29358;
	287: sound1 <=  29297;
	288: sound1 <=  29480;
	289: sound1 <=  29297;
	290: sound1 <=  29724;
	291: sound1 <=  29602;
	292: sound1 <=  29480;
	293: sound1 <=  29236;
	294: sound1 <=  29114;
	295: sound1 <=  29266;
	296: sound1 <=  28992;
	297: sound1 <=  29358;
	298: sound1 <=  29205;
	299: sound1 <=  29266;
	300: sound1 <=  29297;
	301: sound1 <=  29388;
	302: sound1 <=  28809;
	303: sound1 <=  29327;
	304: sound1 <=  29541;
	305: sound1 <=  29205;
	306: sound1 <=  29175;
	307: sound1 <=  29297;
	308: sound1 <=  29266;
	309: sound1 <=  28992;
	310: sound1 <=  29022;
	311: sound1 <=  28809;
	312: sound1 <=  28931;
	313: sound1 <=  28809;
	314: sound1 <=  29083;
	315: sound1 <=  28870;
	316: sound1 <=  28778;
	317: sound1 <=  29114;
	318: sound1 <=  28809;
	319: sound1 <=  28992;
	320: sound1 <=  29236;
	321: sound1 <=  28900;
	322: sound1 <=  28778;
	323: sound1 <=  28748;
	324: sound1 <=  28992;
	325: sound1 <=  28503;
	326: sound1 <=  28595;
	327: sound1 <=  28931;
	328: sound1 <=  28778;
	329: sound1 <=  28717;
	330: sound1 <=  28748;
	331: sound1 <=  28503;
	332: sound1 <=  28137;
	333: sound1 <=  28168;
	334: sound1 <=  28259;
	335: sound1 <=  28412;
	336: sound1 <=  28381;
	337: sound1 <=  28412;
	338: sound1 <=  28778;
	339: sound1 <=  28534;
	340: sound1 <=  28748;
	341: sound1 <=  28992;
	342: sound1 <=  28503;
	343: sound1 <=  28595;
	344: sound1 <=  29175;
	345: sound1 <=  28961;
	346: sound1 <=  28717;
	347: sound1 <=  29083;
	348: sound1 <=  28778;
	349: sound1 <=  28717;
	350: sound1 <=  28625;
	351: sound1 <=  28961;
	352: sound1 <=  29022;
	353: sound1 <=  28656;
	354: sound1 <=  28839;
	355: sound1 <=  29175;
	356: sound1 <=  28809;
	357: sound1 <=  29236;
	358: sound1 <=  29297;
	359: sound1 <=  29327;
	360: sound1 <=  29327;
	361: sound1 <=  29572;
	362: sound1 <=  29633;
	363: sound1 <=  29327;
	364: sound1 <=  29144;
	365: sound1 <=  29419;
	366: sound1 <=  29510;
	367: sound1 <=  29907;
	368: sound1 <=  29388;
	369: sound1 <=  29327;
	370: sound1 <=  29327;
	371: sound1 <=  29175;
	372: sound1 <=  29816;
	373: sound1 <=  29419;
	374: sound1 <=  29388;
	375: sound1 <=  29785;
	376: sound1 <=  29419;
	377: sound1 <=  29297;
	378: sound1 <=  29510;
	379: sound1 <=  29724;
	380: sound1 <=  29449;
	381: sound1 <=  29755;
	382: sound1 <=  29388;
	383: sound1 <=  29266;
	384: sound1 <=  29724;
	385: sound1 <=  29388;
	386: sound1 <=  29388;
	387: sound1 <=  29510;
	388: sound1 <=  29388;
	389: sound1 <=  29114;
	390: sound1 <=  29572;
	391: sound1 <=  28961;
	392: sound1 <=  29449;
	393: sound1 <=  29541;
	394: sound1 <=  29724;
	395: sound1 <=  29327;
	396: sound1 <=  29602;
	397: sound1 <=  29236;
	398: sound1 <=  28961;
	399: sound1 <=  29053;
	400: sound1 <=  29327;
	401: sound1 <=  29205;
	402: sound1 <=  28870;
	403: sound1 <=  29449;
	404: sound1 <=  29419;
	405: sound1 <=  28961;
	406: sound1 <=  29327;
	407: sound1 <=  29266;
	408: sound1 <=  29144;
	409: sound1 <=  29572;
	410: sound1 <=  29480;
	411: sound1 <=  29205;
	412: sound1 <=  29388;
	413: sound1 <=  29724;
	414: sound1 <=  29572;
	415: sound1 <=  29297;
	416: sound1 <=  29480;
	417: sound1 <=  29633;
	418: sound1 <=  30090;
	419: sound1 <=  29846;
	420: sound1 <=  30243;
	421: sound1 <=  30121;
	422: sound1 <=  30090;
	423: sound1 <=  30579;
	424: sound1 <=  30457;
	425: sound1 <=  31189;
	426: sound1 <=  31006;
	427: sound1 <=  31281;
	428: sound1 <=  31006;
	429: sound1 <=  31494;
	430: sound1 <=  32227;
	431: sound1 <=  32440;
	432: sound1 <=  31921;
	433: sound1 <=  31921;
	434: sound1 <=  32104;
	435: sound1 <=  32440;
	436: sound1 <=  32806;
	437: sound1 <=  32562;
	438: sound1 <=  32623;
	439: sound1 <=  32867;
	440: sound1 <=  32501;
	441: sound1 <=  32715;
	442: sound1 <=  33234;
	443: sound1 <=  33112;
	444: sound1 <=  33234;
	445: sound1 <=  33630;
	446: sound1 <=  33813;
	447: sound1 <=  33844;
	448: sound1 <=  34058;
	449: sound1 <=  34058;
	450: sound1 <=  33875;
	451: sound1 <=  34271;
	452: sound1 <=  34210;
	453: sound1 <=  34698;
	454: sound1 <=  34637;
	455: sound1 <=  34729;
	456: sound1 <=  34058;
	457: sound1 <=  35034;
	458: sound1 <=  34973;
	459: sound1 <=  34424;
	460: sound1 <=  34241;
	461: sound1 <=  34637;
	462: sound1 <=  34424;
	463: sound1 <=  34363;
	464: sound1 <=  34119;
	465: sound1 <=  33752;
	466: sound1 <=  34027;
	467: sound1 <=  34027;
	468: sound1 <=  33447;
	469: sound1 <=  33417;
	470: sound1 <=  33173;
	471: sound1 <=  33325;
	472: sound1 <=  32806;
	473: sound1 <=  32562;
	474: sound1 <=  32990;
	475: sound1 <=  32776;
	476: sound1 <=  32135;
	477: sound1 <=  31921;
	478: sound1 <=  31494;
	479: sound1 <=  31067;
	480: sound1 <=  30823;
	481: sound1 <=  31067;
	482: sound1 <=  30182;
	483: sound1 <=  29907;
	484: sound1 <=  30121;
	485: sound1 <=  29449;
	486: sound1 <=  29144;
	487: sound1 <=  28870;
	488: sound1 <=  28442;
	489: sound1 <=  28168;
	490: sound1 <=  28076;
	491: sound1 <=  27527;
	492: sound1 <=  27252;
	493: sound1 <=  27283;
	494: sound1 <=  26733;
	495: sound1 <=  26337;
	496: sound1 <=  26611;
	497: sound1 <=  26154;
	498: sound1 <=  25421;
	499: sound1 <=  25116;
	500: sound1 <=  25055;
	501: sound1 <=  25208;
	502: sound1 <=  24506;
	503: sound1 <=  24353;
	504: sound1 <=  24139;
	505: sound1 <=  24475;
	506: sound1 <=  24445;
	507: sound1 <=  23926;
	508: sound1 <=  24078;
	509: sound1 <=  23987;
	510: sound1 <=  23560;
	511: sound1 <=  23712;
	512: sound1 <=  23956;
	513: sound1 <=  23895;
	514: sound1 <=  23804;
	515: sound1 <=  23773;
	516: sound1 <=  24109;
	517: sound1 <=  23956;
	518: sound1 <=  23529;
	519: sound1 <=  24048;
	520: sound1 <=  24414;
	521: sound1 <=  24963;
	522: sound1 <=  25116;
	523: sound1 <=  24689;
	524: sound1 <=  24780;
	525: sound1 <=  25360;
	526: sound1 <=  25391;
	527: sound1 <=  25177;
	528: sound1 <=  25055;
	529: sound1 <=  25848;
	530: sound1 <=  26093;
	531: sound1 <=  25848;
	532: sound1 <=  26154;
	533: sound1 <=  26245;
	534: sound1 <=  26703;
	535: sound1 <=  27039;
	536: sound1 <=  26611;
	537: sound1 <=  26825;
	538: sound1 <=  27588;
	539: sound1 <=  27344;
	540: sound1 <=  27405;
	541: sound1 <=  27527;
	542: sound1 <=  27557;
	543: sound1 <=  28015;
	544: sound1 <=  28137;
	545: sound1 <=  28320;
	546: sound1 <=  28625;
	547: sound1 <=  27863;
	548: sound1 <=  28687;
	549: sound1 <=  28442;
	550: sound1 <=  28320;
	551: sound1 <=  28412;
	552: sound1 <=  28259;
	553: sound1 <=  28381;
	554: sound1 <=  27985;
	555: sound1 <=  28381;
	556: sound1 <=  28503;
	557: sound1 <=  27924;
	558: sound1 <=  27527;
	559: sound1 <=  27771;
	560: sound1 <=  27893;
	561: sound1 <=  27405;
	562: sound1 <=  27649;
	563: sound1 <=  27039;
	564: sound1 <=  26733;
	565: sound1 <=  26794;
	566: sound1 <=  26459;
	567: sound1 <=  26337;
	568: sound1 <=  26031;
	569: sound1 <=  25726;
	570: sound1 <=  25238;
	571: sound1 <=  24933;
	572: sound1 <=  24872;
	573: sound1 <=  24292;
	574: sound1 <=  23346;
	575: sound1 <=  23346;
	576: sound1 <=  22095;
	577: sound1 <=  20569;
	578: sound1 <=  16785;
	579: sound1 <=  10223;
	580: sound1 <=  -4211;
	581: sound1 <=  -33264;
	582: sound1 <=  -66345;
	583: sound1 <=  -82001;
	584: sound1 <=  -80841;
	585: sound1 <=  -65796;
	586: sound1 <=  -41351;
	587: sound1 <=  -11658;
	588: sound1 <=  21759;
	589: sound1 <=  54352;
	590: sound1 <=  83435;
	591: sound1 <=  108490;
	592: sound1 <=  128571;
	593: sound1 <=  145996;
	594: sound1 <=  160767;
	595: sound1 <=  173553;
	596: sound1 <=  184113;
	597: sound1 <=  193146;
	598: sound1 <=  200714;
	599: sound1 <=  205536;
	600: sound1 <=  208862;
	601: sound1 <=  209351;
	602: sound1 <=  207611;
	603: sound1 <=  201813;
	604: sound1 <=  193237;
	605: sound1 <=  182007;
	606: sound1 <=  167816;
	607: sound1 <=  151245;
	608: sound1 <=  132751;
	609: sound1 <=  112457;
	610: sound1 <=  90820;
	611: sound1 <=  67139;
	612: sound1 <=  42236;
	613: sound1 <=  17212;
	614: sound1 <=  -9460;
	615: sound1 <=  -35217;
	616: sound1 <=  -61676;
	617: sound1 <=  -88562;
	618: sound1 <=  -117035;
	619: sound1 <=  -145721;
	620: sound1 <=  -175995;
	621: sound1 <=  -204926;
	622: sound1 <=  -234039;
	623: sound1 <=  -261993;
	624: sound1 <=  -279205;
	625: sound1 <=  -283051;
	626: sound1 <=  -280212;
	627: sound1 <=  -276367;
	628: sound1 <=  -271942;
	629: sound1 <=  -266174;
	630: sound1 <=  -260284;
	631: sound1 <=  -253967;
	632: sound1 <=  -244110;
	633: sound1 <=  -232025;
	634: sound1 <=  -220306;
	635: sound1 <=  -212982;
	636: sound1 <=  -208191;
	637: sound1 <=  -204620;
	638: sound1 <=  -201569;
	639: sound1 <=  -198425;
	640: sound1 <=  -194366;
	641: sound1 <=  -188293;
	642: sound1 <=  -180847;
	643: sound1 <=  -171661;
	644: sound1 <=  -161743;
	645: sound1 <=  -150452;
	646: sound1 <=  -137848;
	647: sound1 <=  -124237;
	648: sound1 <=  -109253;
	649: sound1 <=  -91278;
	650: sound1 <=  -67108;
	651: sound1 <=  -35675;
	652: sound1 <=  732;
	653: sound1 <=  39795;
	654: sound1 <=  81055;
	655: sound1 <=  121155;
	656: sound1 <=  157776;
	657: sound1 <=  183777;
	658: sound1 <=  196014;
	659: sound1 <=  191467;
	660: sound1 <=  168274;
	661: sound1 <=  123962;
	662: sound1 <=  54962;
	663: sound1 <=  -29846;
	664: sound1 <=  -73395;
	665: sound1 <=  -75256;
	666: sound1 <=  -73486;
	667: sound1 <=  -67688;
	668: sound1 <=  -60577;
	669: sound1 <=  -53192;
	670: sound1 <=  -43518;
	671: sound1 <=  -32959;
	672: sound1 <=  -21484;
	673: sound1 <=  -8484;
	674: sound1 <=  7965;
	675: sound1 <=  25208;
	676: sound1 <=  70435;
	677: sound1 <=  171570;
	678: sound1 <=  313873;
	679: sound1 <=  421356;
	680: sound1 <=  493469;
	681: sound1 <=  556213;
	682: sound1 <=  447418;
	683: sound1 <=  333954;
	684: sound1 <=  344086;
	685: sound1 <=  351227;
	686: sound1 <=  366119;
	687: sound1 <=  376129;
	688: sound1 <=  385681;
	689: sound1 <=  392609;
	690: sound1 <=  397278;
	691: sound1 <=  399048;
	692: sound1 <=  399963;
	693: sound1 <=  398376;
	694: sound1 <=  394073;
	695: sound1 <=  389221;
	696: sound1 <=  382263;
	697: sound1 <=  374451;
	698: sound1 <=  365936;
	699: sound1 <=  356842;
	700: sound1 <=  348053;
	701: sound1 <=  340118;
	702: sound1 <=  337585;
	703: sound1 <=  363770;
	704: sound1 <=  367676;
	705: sound1 <=  297882;
	706: sound1 <=  167725;
	707: sound1 <=  25543;
	708: sound1 <=  -106598;
	709: sound1 <=  -167908;
	710: sound1 <=  -178131;
	711: sound1 <=  -184662;
	712: sound1 <=  -185059;
	713: sound1 <=  -182373;
	714: sound1 <=  -174774;
	715: sound1 <=  -169220;
	716: sound1 <=  -175293;
	717: sound1 <=  -185089;
	718: sound1 <=  -192810;
	719: sound1 <=  -198364;
	720: sound1 <=  -201630;
	721: sound1 <=  -201782;
	722: sound1 <=  -200623;
	723: sound1 <=  -197632;
	724: sound1 <=  -192780;
	725: sound1 <=  -187347;
	726: sound1 <=  -181610;
	727: sound1 <=  -176300;
	728: sound1 <=  -178711;
	729: sound1 <=  -190613;
	730: sound1 <=  -204712;
	731: sound1 <=  -205017;
	732: sound1 <=  -202881;
	733: sound1 <=  -184448;
	734: sound1 <=  -135376;
	735: sound1 <=  -105194;
	736: sound1 <=  -95398;
	737: sound1 <=  -93567;
	738: sound1 <=  -99060;
	739: sound1 <=  -104553;
	740: sound1 <=  -107727;
	741: sound1 <=  -109131;
	742: sound1 <=  -107819;
	743: sound1 <=  -103607;
	744: sound1 <=  -96588;
	745: sound1 <=  -83954;
	746: sound1 <=  -61646;
	747: sound1 <=  -21210;
	748: sound1 <=  22003;
	749: sound1 <=  51788;
	750: sound1 <=  75562;
	751: sound1 <=  96527;
	752: sound1 <=  122711;
	753: sound1 <=  157501;
	754: sound1 <=  195038;
	755: sound1 <=  236328;
	756: sound1 <=  286163;
	757: sound1 <=  339142;
	758: sound1 <=  400818;
	759: sound1 <=  464783;
	760: sound1 <=  518585;
	761: sound1 <=  546661;
	762: sound1 <=  550873;
	763: sound1 <=  534058;
	764: sound1 <=  489777;
	765: sound1 <=  424072;
	766: sound1 <=  366241;
	767: sound1 <=  338989;
	768: sound1 <=  341980;
	769: sound1 <=  360260;
	770: sound1 <=  383301;
	771: sound1 <=  401794;
	772: sound1 <=  412292;
	773: sound1 <=  421448;
	774: sound1 <=  429504;
	775: sound1 <=  427460;
	776: sound1 <=  419312;
	777: sound1 <=  408356;
	778: sound1 <=  394196;
	779: sound1 <=  369843;
	780: sound1 <=  337067;
	781: sound1 <=  263580;
	782: sound1 <=  140259;
	783: sound1 <=  42542;
	784: sound1 <=  -22675;
	785: sound1 <=  -62012;
	786: sound1 <=  -78766;
	787: sound1 <=  -80414;
	788: sound1 <=  -73181;
	789: sound1 <=  -58655;
	790: sound1 <=  -44678;
	791: sound1 <=  -36621;
	792: sound1 <=  -28625;
	793: sound1 <=  -22461;
	794: sound1 <=  -24475;
	795: sound1 <=  -37842;
	796: sound1 <=  -55573;
	797: sound1 <=  -77728;
	798: sound1 <=  -102478;
	799: sound1 <=  -120544;
	800: sound1 <=  -124146;
	801: sound1 <=  -115479;
	802: sound1 <=  -100708;
	803: sound1 <=  -82001;
	804: sound1 <=  -49957;
	805: sound1 <=  3448;
	806: sound1 <=  79803;
	807: sound1 <=  162018;
	808: sound1 <=  227905;
	809: sound1 <=  260590;
	810: sound1 <=  277679;
	811: sound1 <=  277313;
	812: sound1 <=  263000;
	813: sound1 <=  249054;
	814: sound1 <=  236969;
	815: sound1 <=  227722;
	816: sound1 <=  222290;
	817: sound1 <=  214478;
	818: sound1 <=  199310;
	819: sound1 <=  166565;
	820: sound1 <=  67230;
	821: sound1 <=  -251709;
	822: sound1 <=  -504456;
	823: sound1 <=  -524506;
	824: sound1 <=  -542206;
	825: sound1 <=  -545227;
	826: sound1 <=  -546173;
	827: sound1 <=  -540741;
	828: sound1 <=  -532715;
	829: sound1 <=  -518066;
	830: sound1 <=  -491516;
	831: sound1 <=  -443024;
	832: sound1 <=  -306122;
	833: sound1 <=  -130463;
	834: sound1 <=  -4639;
	835: sound1 <=  72968;
	836: sound1 <=  146790;
	837: sound1 <=  220459;
	838: sound1 <=  285645;
	839: sound1 <=  326355;
	840: sound1 <=  322601;
	841: sound1 <=  296722;
	842: sound1 <=  270264;
	843: sound1 <=  163361;
	844: sound1 <=  -34149;
	845: sound1 <=  -147736;
	846: sound1 <=  -177551;
	847: sound1 <=  -142487;
	848: sound1 <=  -83923;
	849: sound1 <=  -43488;
	850: sound1 <=  -14740;
	851: sound1 <=  -11261;
	852: sound1 <=  -73242;
	853: sound1 <=  -344788;
	854: sound1 <=  -477051;
	855: sound1 <=  -470032;
	856: sound1 <=  -494446;
	857: sound1 <=  -501556;
	858: sound1 <=  -518097;
	859: sound1 <=  -525726;
	860: sound1 <=  -526459;
	861: sound1 <=  -512665;
	862: sound1 <=  -499878;
	863: sound1 <=  -481934;
	864: sound1 <=  -464386;
	865: sound1 <=  -443176;
	866: sound1 <=  -418915;
	867: sound1 <=  -356140;
	868: sound1 <=  -214935;
	869: sound1 <=  -87524;
	870: sound1 <=  22034;
	871: sound1 <=  105072;
	872: sound1 <=  227600;
	873: sound1 <=  377960;
	874: sound1 <=  472290;
	875: sound1 <=  499542;
	876: sound1 <=  485291;
	877: sound1 <=  466614;
	878: sound1 <=  447205;
	879: sound1 <=  427216;
	880: sound1 <=  407410;
	881: sound1 <=  385254;
	882: sound1 <=  362274;
	883: sound1 <=  332672;
	884: sound1 <=  291199;
	885: sound1 <=  252380;
	886: sound1 <=  230591;
	887: sound1 <=  205841;
	888: sound1 <=  168091;
	889: sound1 <=  -26215;
	890: sound1 <=  -254486;
	891: sound1 <=  -369568;
	892: sound1 <=  -412445;
	893: sound1 <=  -398224;
	894: sound1 <=  -375275;
	895: sound1 <=  -325439;
	896: sound1 <=  -273010;
	897: sound1 <=  -241943;
	898: sound1 <=  -231506;
	899: sound1 <=  -232239;
	900: sound1 <=  -222534;
	901: sound1 <=  -201874;
	902: sound1 <=  -178436;
	903: sound1 <=  -146729;
	904: sound1 <=  -97534;
	905: sound1 <=  -24170;
	906: sound1 <=  -49805;
	907: sound1 <=  -191071;
	908: sound1 <=  -221191;
	909: sound1 <=  -236633;
	910: sound1 <=  -249329;
	911: sound1 <=  -257538;
	912: sound1 <=  -263245;
	913: sound1 <=  -265625;
	914: sound1 <=  -266724;
	915: sound1 <=  -258575;
	916: sound1 <=  -248291;
	917: sound1 <=  -237640;
	918: sound1 <=  -219604;
	919: sound1 <=  -210846;
	920: sound1 <=  -214142;
	921: sound1 <=  -214203;
	922: sound1 <=  -206909;
	923: sound1 <=  -205780;
	924: sound1 <=  -205017;
	925: sound1 <=  -147217;
	926: sound1 <=  -28625;
	927: sound1 <=  80078;
	928: sound1 <=  183655;
	929: sound1 <=  262360;
	930: sound1 <=  332458;
	931: sound1 <=  411163;
	932: sound1 <=  484894;
	933: sound1 <=  553345;
	934: sound1 <=  593262;
	935: sound1 <=  588226;
	936: sound1 <=  578949;
	937: sound1 <=  567169;
	938: sound1 <=  553680;
	939: sound1 <=  537201;
	940: sound1 <=  533417;
	941: sound1 <=  557068;
	942: sound1 <=  566742;
	943: sound1 <=  556976;
	944: sound1 <=  536346;
	945: sound1 <=  509460;
	946: sound1 <=  474579;
	947: sound1 <=  433289;
	948: sound1 <=  394226;
	949: sound1 <=  359039;
	950: sound1 <=  333771;
	951: sound1 <=  316772;
	952: sound1 <=  298859;
	953: sound1 <=  280243;
	954: sound1 <=  264618;
	955: sound1 <=  247406;
	956: sound1 <=  231537;
	957: sound1 <=  215179;
	958: sound1 <=  217346;
	959: sound1 <=  219788;
	960: sound1 <=  196136;
	961: sound1 <=  167908;
	962: sound1 <=  128326;
	963: sound1 <=  80261;
	964: sound1 <=  18494;
	965: sound1 <=  -41290;
	966: sound1 <=  -106628;
	967: sound1 <=  -159821;
	968: sound1 <=  -291412;
	969: sound1 <=  -419342;
	970: sound1 <=  -427032;
	971: sound1 <=  -455627;
	972: sound1 <=  -473877;
	973: sound1 <=  -486450;
	974: sound1 <=  -490051;
	975: sound1 <=  -491791;
	976: sound1 <=  -484985;
	977: sound1 <=  -482147;
	978: sound1 <=  -474976;
	979: sound1 <=  -469238;
	980: sound1 <=  -457703;
	981: sound1 <=  -455688;
	982: sound1 <=  -457031;
	983: sound1 <=  -450653;
	984: sound1 <=  -427399;
	985: sound1 <=  -398834;
	986: sound1 <=  -303070;
	987: sound1 <=  -298248;
	988: sound1 <=  -313171;
	989: sound1 <=  -247162;
	990: sound1 <=  -163788;
	991: sound1 <=  -76599;
	992: sound1 <=  23682;
	993: sound1 <=  -24750;
	994: sound1 <=  -195953;
	995: sound1 <=  -108704;
	996: sound1 <=  -10620;
	997: sound1 <=  -30304;
	998: sound1 <=  -191925;
	999: sound1 <=  -175598;
	1000: sound1 <=  -123566;
	1001: sound1 <=  -45563;
	1002: sound1 <=  -105865;
	1003: sound1 <=  -144623;
	1004: sound1 <=  -130127;
	1005: sound1 <=  -123352;
	1006: sound1 <=  -110901;
	1007: sound1 <=  -141724;
	1008: sound1 <=  -133759;
	1009: sound1 <=  -98969;
	1010: sound1 <=  -21423;
	1011: sound1 <=  79193;
	1012: sound1 <=  488;
	1013: sound1 <=  -19165;
	1014: sound1 <=  6744;
	1015: sound1 <=  44800;
	1016: sound1 <=  137909;
	1017: sound1 <=  239136;
	1018: sound1 <=  341248;
	1019: sound1 <=  425690;
	1020: sound1 <=  496490;
	1021: sound1 <=  526947;
	1022: sound1 <=  559479;
	1023: sound1 <=  468597;
	1024: sound1 <=  88348;
	1025: sound1 <=  24414;
	1026: sound1 <=  24841;
	1027: sound1 <=  23712;
	1028: sound1 <=  33142;
	1029: sound1 <=  49591;
	1030: sound1 <=  72266;
	1031: sound1 <=  108643;
	1032: sound1 <=  155304;
	1033: sound1 <=  237091;
	1034: sound1 <=  394409;
	1035: sound1 <=  507202;
	1036: sound1 <=  579956;
	1037: sound1 <=  654266;
	1038: sound1 <=  660370;
	1039: sound1 <=  711914;
	1040: sound1 <=  721802;
	1041: sound1 <=  685272;
	1042: sound1 <=  665253;
	1043: sound1 <=  649628;
	1044: sound1 <=  625946;
	1045: sound1 <=  644592;
	1046: sound1 <=  644897;
	1047: sound1 <=  602417;
	1048: sound1 <=  565552;
	1049: sound1 <=  575592;
	1050: sound1 <=  579926;
	1051: sound1 <=  549042;
	1052: sound1 <=  517517;
	1053: sound1 <=  496399;
	1054: sound1 <=  501007;
	1055: sound1 <=  483856;
	1056: sound1 <=  459503;
	1057: sound1 <=  440094;
	1058: sound1 <=  426208;
	1059: sound1 <=  421021;
	1060: sound1 <=  390808;
	1061: sound1 <=  331757;
	1062: sound1 <=  245087;
	1063: sound1 <=  220825;
	1064: sound1 <=  267059;
	1065: sound1 <=  258972;
	1066: sound1 <=  260284;
	1067: sound1 <=  249786;
	1068: sound1 <=  237061;
	1069: sound1 <=  218506;
	1070: sound1 <=  174255;
	1071: sound1 <=  118103;
	1072: sound1 <=  72357;
	1073: sound1 <=  28259;
	1074: sound1 <=  -42480;
	1075: sound1 <=  3723;
	1076: sound1 <=  3937;
	1077: sound1 <=  -39764;
	1078: sound1 <=  -65979;
	1079: sound1 <=  -100403;
	1080: sound1 <=  -143646;
	1081: sound1 <=  -281036;
	1082: sound1 <=  -333405;
	1083: sound1 <=  -369415;
	1084: sound1 <=  -411194;
	1085: sound1 <=  -457825;
	1086: sound1 <=  -481842;
	1087: sound1 <=  -473267;
	1088: sound1 <=  -462799;
	1089: sound1 <=  -460663;
	1090: sound1 <=  -455139;
	1091: sound1 <=  -452301;
	1092: sound1 <=  -438568;
	1093: sound1 <=  -420746;
	1094: sound1 <=  -422180;
	1095: sound1 <=  -415253;
	1096: sound1 <=  -379639;
	1097: sound1 <=  -312317;
	1098: sound1 <=  -235565;
	1099: sound1 <=  -185638;
	1100: sound1 <=  -74554;
	1101: sound1 <=  -8728;
	1102: sound1 <=  35950;
	1103: sound1 <=  67841;
	1104: sound1 <=  108032;
	1105: sound1 <=  130737;
	1106: sound1 <=  168945;
	1107: sound1 <=  64209;
	1108: sound1 <=  -340668;
	1109: sound1 <=  -366699;
	1110: sound1 <=  -365692;
	1111: sound1 <=  -370087;
	1112: sound1 <=  -348694;
	1113: sound1 <=  -316589;
	1114: sound1 <=  -284088;
	1115: sound1 <=  -210358;
	1116: sound1 <=  -112518;
	1117: sound1 <=  -61310;
	1118: sound1 <=  20721;
	1119: sound1 <=  -188934;
	1120: sound1 <=  -342285;
	1121: sound1 <=  -320221;
	1122: sound1 <=  -317413;
	1123: sound1 <=  -272827;
	1124: sound1 <=  -202057;
	1125: sound1 <=  -84534;
	1126: sound1 <=  -22980;
	1127: sound1 <=  22308;
	1128: sound1 <=  65308;
	1129: sound1 <=  81879;
	1130: sound1 <=  35065;
	1131: sound1 <=  -29999;
	1132: sound1 <=  2747;
	1133: sound1 <=  24384;
	1134: sound1 <=  -27740;
	1135: sound1 <=  -85724;
	1136: sound1 <=  -133301;
	1137: sound1 <=  -164520;
	1138: sound1 <=  -164032;
	1139: sound1 <=  -141235;
	1140: sound1 <=  -127960;
	1141: sound1 <=  -124298;
	1142: sound1 <=  -130951;
	1143: sound1 <=  -131531;
	1144: sound1 <=  -132660;
	1145: sound1 <=  -122772;
	1146: sound1 <=  -103455;
	1147: sound1 <=  -90057;
	1148: sound1 <=  -53741;
	1149: sound1 <=  67047;
	1150: sound1 <=  189301;
	1151: sound1 <=  223419;
	1152: sound1 <=  235229;
	1153: sound1 <=  231934;
	1154: sound1 <=  254944;
	1155: sound1 <=  131714;
	1156: sound1 <=  -259674;
	1157: sound1 <=  -258331;
	1158: sound1 <=  -246460;
	1159: sound1 <=  -186066;
	1160: sound1 <=  -147980;
	1161: sound1 <=  -162384;
	1162: sound1 <=  -152954;
	1163: sound1 <=  -146362;
	1164: sound1 <=  -137451;
	1165: sound1 <=  -130219;
	1166: sound1 <=  -118225;
	1167: sound1 <=  -95581;
	1168: sound1 <=  -58685;
	1169: sound1 <=  -2045;
	1170: sound1 <=  110870;
	1171: sound1 <=  292053;
	1172: sound1 <=  423370;
	1173: sound1 <=  491852;
	1174: sound1 <=  560944;
	1175: sound1 <=  636810;
	1176: sound1 <=  692719;
	1177: sound1 <=  712585;
	1178: sound1 <=  675812;
	1179: sound1 <=  601868;
	1180: sound1 <=  486877;
	1181: sound1 <=  341614;
	1182: sound1 <=  276489;
	1183: sound1 <=  282379;
	1184: sound1 <=  278870;
	1185: sound1 <=  279938;
	1186: sound1 <=  272369;
	1187: sound1 <=  281403;
	1188: sound1 <=  291718;
	1189: sound1 <=  289001;
	1190: sound1 <=  279541;
	1191: sound1 <=  251831;
	1192: sound1 <=  225647;
	1193: sound1 <=  232178;
	1194: sound1 <=  255524;
	1195: sound1 <=  285553;
	1196: sound1 <=  306671;
	1197: sound1 <=  326355;
	1198: sound1 <=  343170;
	1199: sound1 <=  332550;
	1200: sound1 <=  312775;
	1201: sound1 <=  268982;
	1202: sound1 <=  209991;
	1203: sound1 <=  156372;
	1204: sound1 <=  70374;
	1205: sound1 <=  -25146;
	1206: sound1 <=  -113220;
	1207: sound1 <=  -111511;
	1208: sound1 <=  -118652;
	1209: sound1 <=  -177917;
	1210: sound1 <=  -221191;
	1211: sound1 <=  -238525;
	1212: sound1 <=  -244263;
	1213: sound1 <=  -256195;
	1214: sound1 <=  -269501;
	1215: sound1 <=  -282654;
	1216: sound1 <=  -287415;
	1217: sound1 <=  -294403;
	1218: sound1 <=  -309418;
	1219: sound1 <=  -315460;
	1220: sound1 <=  -309540;
	1221: sound1 <=  -308044;
	1222: sound1 <=  -325623;
	1223: sound1 <=  -357605;
	1224: sound1 <=  -378693;
	1225: sound1 <=  -373505;
	1226: sound1 <=  -364166;
	1227: sound1 <=  -367706;
	1228: sound1 <=  -392151;
	1229: sound1 <=  -404816;
	1230: sound1 <=  -383789;
	1231: sound1 <=  -341644;
	1232: sound1 <=  -273804;
	1233: sound1 <=  -203766;
	1234: sound1 <=  -173431;
	1235: sound1 <=  -192596;
	1236: sound1 <=  -188324;
	1237: sound1 <=  -171997;
	1238: sound1 <=  -154205;
	1239: sound1 <=  -192749;
	1240: sound1 <=  -206329;
	1241: sound1 <=  -205719;
	1242: sound1 <=  -194672;
	1243: sound1 <=  -173157;
	1244: sound1 <=  -165192;
	1245: sound1 <=  -147797;
	1246: sound1 <=  -136292;
	1247: sound1 <=  -121735;
	1248: sound1 <=  -123932;
	1249: sound1 <=  -121002;
	1250: sound1 <=  -90271;
	1251: sound1 <=  -69397;
	1252: sound1 <=  -5493;
	1253: sound1 <=  22095;
	1254: sound1 <=  43579;
	1255: sound1 <=  104370;
	1256: sound1 <=  153259;
	1257: sound1 <=  225647;
	1258: sound1 <=  286469;
	1259: sound1 <=  337311;
	1260: sound1 <=  375458;
	1261: sound1 <=  405975;
	1262: sound1 <=  391693;
	1263: sound1 <=  369171;
	1264: sound1 <=  344727;
	1265: sound1 <=  280457;
	1266: sound1 <=  233978;
	1267: sound1 <=  227234;
	1268: sound1 <=  191559;
	1269: sound1 <=  170776;
	1270: sound1 <=  170013;
	1271: sound1 <=  179932;
	1272: sound1 <=  176666;
	1273: sound1 <=  163940;
	1274: sound1 <=  166779;
	1275: sound1 <=  200958;
	1276: sound1 <=  240356;
	1277: sound1 <=  256989;
	1278: sound1 <=  281158;
	1279: sound1 <=  303558;
	1280: sound1 <=  288116;
	1281: sound1 <=  267914;
	1282: sound1 <=  213684;
	1283: sound1 <=  139008;
	1284: sound1 <=  56763;
	1285: sound1 <=  -42480;
	1286: sound1 <=  -49988;
	1287: sound1 <=  -74738;
	1288: sound1 <=  -83649;
	1289: sound1 <=  -82886;
	1290: sound1 <=  -80627;
	1291: sound1 <=  -76965;
	1292: sound1 <=  -84198;
	1293: sound1 <=  -108032;
	1294: sound1 <=  -124268;
	1295: sound1 <=  -120697;
	1296: sound1 <=  -123840;
	1297: sound1 <=  -138428;
	1298: sound1 <=  -135010;
	1299: sound1 <=  -118927;
	1300: sound1 <=  -109406;
	1301: sound1 <=  -129913;
	1302: sound1 <=  -126831;
	1303: sound1 <=  -73578;
	1304: sound1 <=  33447;
	1305: sound1 <=  133514;
	1306: sound1 <=  204498;
	1307: sound1 <=  308075;
	1308: sound1 <=  391479;
	1309: sound1 <=  467773;
	1310: sound1 <=  554047;
	1311: sound1 <=  616119;
	1312: sound1 <=  638458;
	1313: sound1 <=  592834;
	1314: sound1 <=  549072;
	1315: sound1 <=  527588;
	1316: sound1 <=  525269;
	1317: sound1 <=  534515;
	1318: sound1 <=  541290;
	1319: sound1 <=  531433;
	1320: sound1 <=  514069;
	1321: sound1 <=  518463;
	1322: sound1 <=  507996;
	1323: sound1 <=  464355;
	1324: sound1 <=  425537;
	1325: sound1 <=  406616;
	1326: sound1 <=  373596;
	1327: sound1 <=  350189;
	1328: sound1 <=  334564;
	1329: sound1 <=  319366;
	1330: sound1 <=  268585;
	1331: sound1 <=  221191;
	1332: sound1 <=  197540;
	1333: sound1 <=  182648;
	1334: sound1 <=  199493;
	1335: sound1 <=  202148;
	1336: sound1 <=  183105;
	1337: sound1 <=  147186;
	1338: sound1 <=  107910;
	1339: sound1 <=  77484;
	1340: sound1 <=  49194;
	1341: sound1 <=  27435;
	1342: sound1 <=  -26611;
	1343: sound1 <=  -96985;
	1344: sound1 <=  -151245;
	1345: sound1 <=  -205994;
	1346: sound1 <=  -251678;
	1347: sound1 <=  -330933;
	1348: sound1 <=  -353729;
	1349: sound1 <=  -394623;
	1350: sound1 <=  -416443;
	1351: sound1 <=  -419830;
	1352: sound1 <=  -433624;
	1353: sound1 <=  -426819;
	1354: sound1 <=  -405182;
	1355: sound1 <=  -386658;
	1356: sound1 <=  -406891;
	1357: sound1 <=  -386414;
	1358: sound1 <=  -369019;
	1359: sound1 <=  -352814;
	1360: sound1 <=  -334564;
	1361: sound1 <=  -350830;
	1362: sound1 <=  -377167;
	1363: sound1 <=  -399719;
	1364: sound1 <=  -386414;
	1365: sound1 <=  -349274;
	1366: sound1 <=  -282410;
	1367: sound1 <=  -234100;
	1368: sound1 <=  -207520;
	1369: sound1 <=  -186127;
	1370: sound1 <=  -171753;
	1371: sound1 <=  -173340;
	1372: sound1 <=  -178833;
	1373: sound1 <=  -175720;
	1374: sound1 <=  -165924;
	1375: sound1 <=  -163239;
	1376: sound1 <=  -152130;
	1377: sound1 <=  -140686;
	1378: sound1 <=  -128021;
	1379: sound1 <=  -113708;
	1380: sound1 <=  -112213;
	1381: sound1 <=  -104614;
	1382: sound1 <=  -98999;
	1383: sound1 <=  -86487;
	1384: sound1 <=  -56519;
	1385: sound1 <=  -55450;
	1386: sound1 <=  -34424;
	1387: sound1 <=  -81268;
	1388: sound1 <=  -95490;
	1389: sound1 <=  -39886;
	1390: sound1 <=  -47333;
	1391: sound1 <=  104553;
	1392: sound1 <=  54596;
	1393: sound1 <=  215668;
	1394: sound1 <=  246643;
	1395: sound1 <=  143036;
	1396: sound1 <=  248718;
	1397: sound1 <=  260803;
	1398: sound1 <=  317932;
	1399: sound1 <=  375183;
	1400: sound1 <=  433838;
	1401: sound1 <=  319000;
	1402: sound1 <=  126984;
	1403: sound1 <=  133301;
	1404: sound1 <=  125092;
	1405: sound1 <=  151825;
	1406: sound1 <=  144501;
	1407: sound1 <=  135590;
	1408: sound1 <=  173157;
	1409: sound1 <=  256348;
	1410: sound1 <=  315948;
	1411: sound1 <=  340759;
	1412: sound1 <=  395508;
	1413: sound1 <=  427856;
	1414: sound1 <=  371033;
	1415: sound1 <=  384369;
	1416: sound1 <=  480225;
	1417: sound1 <=  504028;
	1418: sound1 <=  488342;
	1419: sound1 <=  418915;
	1420: sound1 <=  353149;
	1421: sound1 <=  317291;
	1422: sound1 <=  299408;
	1423: sound1 <=  298706;
	1424: sound1 <=  315369;
	1425: sound1 <=  329285;
	1426: sound1 <=  331848;
	1427: sound1 <=  321960;
	1428: sound1 <=  310730;
	1429: sound1 <=  172882;
	1430: sound1 <=  71533;
	1431: sound1 <=  -21820;
	1432: sound1 <=  -95673;
	1433: sound1 <=  -164642;
	1434: sound1 <=  -202423;
	1435: sound1 <=  -194397;
	1436: sound1 <=  -170410;
	1437: sound1 <=  -123718;
	1438: sound1 <=  -99121;
	1439: sound1 <=  -74982;
	1440: sound1 <=  -77759;
	1441: sound1 <=  -58563;
	1442: sound1 <=  -23041;
	1443: sound1 <=  24719;
	1444: sound1 <=  94696;
	1445: sound1 <=  121002;
	1446: sound1 <=  149750;
	1447: sound1 <=  167542;
	1448: sound1 <=  176819;
	1449: sound1 <=  192078;
	1450: sound1 <=  196503;
	1451: sound1 <=  184082;
	1452: sound1 <=  180817;
	1453: sound1 <=  213165;
	1454: sound1 <=  199707;
	1455: sound1 <=  133514;
	1456: sound1 <=  106934;
	1457: sound1 <=  89935;
	1458: sound1 <=  51453;
	1459: sound1 <=  45288;
	1460: sound1 <=  -7263;
	1461: sound1 <=  -42633;
	1462: sound1 <=  -91217;
	1463: sound1 <=  -168243;
	1464: sound1 <=  -222321;
	1465: sound1 <=  -250122;
	1466: sound1 <=  -261566;
	1467: sound1 <=  -308258;
	1468: sound1 <=  -359924;
	1469: sound1 <=  -418793;
	1470: sound1 <=  -455627;
	1471: sound1 <=  -485657;
	1472: sound1 <=  -518738;
	1473: sound1 <=  -559692;
	1474: sound1 <=  -559296;
	1475: sound1 <=  -544220;
	1476: sound1 <=  -518768;
	1477: sound1 <=  -506012;
	1478: sound1 <=  -495392;
	1479: sound1 <=  -481781;
	1480: sound1 <=  -452026;
	1481: sound1 <=  -403717;
	1482: sound1 <=  -359528;
	1483: sound1 <=  -323242;
	1484: sound1 <=  -304962;
	1485: sound1 <=  -290253;
	1486: sound1 <=  -270294;
	1487: sound1 <=  -227081;
	1488: sound1 <=  -138306;
	1489: sound1 <=  -17609;
	1490: sound1 <=  82916;
	1491: sound1 <=  160614;
	1492: sound1 <=  235352;
	1493: sound1 <=  317200;
	1494: sound1 <=  347565;
	1495: sound1 <=  361420;
	1496: sound1 <=  354004;
	1497: sound1 <=  368378;
	1498: sound1 <=  385010;
	1499: sound1 <=  385773;
	1500: sound1 <=  384674;
	1501: sound1 <=  374237;
	1502: sound1 <=  349701;
	1503: sound1 <=  325317;
	1504: sound1 <=  326508;
	1505: sound1 <=  319031;
	1506: sound1 <=  287598;
	1507: sound1 <=  268005;
	1508: sound1 <=  291138;
	1509: sound1 <=  304749;
	1510: sound1 <=  282227;
	1511: sound1 <=  243103;
	1512: sound1 <=  230591;
	1513: sound1 <=  213318;
	1514: sound1 <=  207550;
	1515: sound1 <=  199677;
	1516: sound1 <=  184479;
	1517: sound1 <=  161652;
	1518: sound1 <=  106262;
	1519: sound1 <=  88470;
	1520: sound1 <=  86700;
	1521: sound1 <=  45410;
	1522: sound1 <=  19318;
	1523: sound1 <=  8606;
	1524: sound1 <=  -21454;
	1525: sound1 <=  -53528;
	1526: sound1 <=  -97168;
	1527: sound1 <=  -141998;
	1528: sound1 <=  -374786;
	1529: sound1 <=  -456451;
	1530: sound1 <=  -443024;
	1531: sound1 <=  -448242;
	1532: sound1 <=  -429382;
	1533: sound1 <=  -422760;
	1534: sound1 <=  -396271;
	1535: sound1 <=  -369293;
	1536: sound1 <=  -333649;
	1537: sound1 <=  -297333;
	1538: sound1 <=  -291199;
	1539: sound1 <=  -304169;
	1540: sound1 <=  -314789;
	1541: sound1 <=  -305634;
	1542: sound1 <=  -306122;
	1543: sound1 <=  -288391;
	1544: sound1 <=  -282440;
	1545: sound1 <=  -246490;
	1546: sound1 <=  -261993;
	1547: sound1 <=  -290375;
	1548: sound1 <=  -276031;
	1549: sound1 <=  -268738;
	1550: sound1 <=  -240417;
	1551: sound1 <=  -218689;
	1552: sound1 <=  -206329;
	1553: sound1 <=  -216492;
	1554: sound1 <=  -236176;
	1555: sound1 <=  -240509;
	1556: sound1 <=  -227936;
	1557: sound1 <=  -175873;
	1558: sound1 <=  -103943;
	1559: sound1 <=  -28046;
	1560: sound1 <=  23315;
	1561: sound1 <=  91553;
	1562: sound1 <=  156921;
	1563: sound1 <=  207153;
	1564: sound1 <=  260529;
	1565: sound1 <=  313171;
	1566: sound1 <=  314270;
	1567: sound1 <=  298676;
	1568: sound1 <=  292603;
	1569: sound1 <=  299469;
	1570: sound1 <=  322784;
	1571: sound1 <=  337219;
	1572: sound1 <=  325287;
	1573: sound1 <=  315887;
	1574: sound1 <=  304840;
	1575: sound1 <=  308105;
	1576: sound1 <=  311768;
	1577: sound1 <=  295685;
	1578: sound1 <=  280579;
	1579: sound1 <=  290314;
	1580: sound1 <=  338226;
	1581: sound1 <=  332947;
	1582: sound1 <=  304352;
	1583: sound1 <=  292114;
	1584: sound1 <=  297852;
	1585: sound1 <=  313904;
	1586: sound1 <=  319855;
	1587: sound1 <=  286438;
	1588: sound1 <=  257202;
	1589: sound1 <=  196716;
	1590: sound1 <=  166687;
	1591: sound1 <=  -4181;
	1592: sound1 <=  -315460;
	1593: sound1 <=  -341461;
	1594: sound1 <=  -334351;
	1595: sound1 <=  -285187;
	1596: sound1 <=  -237213;
	1597: sound1 <=  -195282;
	1598: sound1 <=  -153290;
	1599: sound1 <=  -118774;
	1600: sound1 <=  -95276;
	1601: sound1 <=  -99152;
	1602: sound1 <=  -106293;
	1603: sound1 <=  -105530;
	1604: sound1 <=  -94360;
	1605: sound1 <=  -55817;
	1606: sound1 <=  -11139;
	1607: sound1 <=  74677;
	1608: sound1 <=  131226;
	1609: sound1 <=  194000;
	1610: sound1 <=  252167;
	1611: sound1 <=  279022;
	1612: sound1 <=  309692;
	1613: sound1 <=  350952;
	1614: sound1 <=  392609;
	1615: sound1 <=  441376;
	1616: sound1 <=  441437;
	1617: sound1 <=  423889;
	1618: sound1 <=  427643;
	1619: sound1 <=  445007;
	1620: sound1 <=  463257;
	1621: sound1 <=  465485;
	1622: sound1 <=  449982;
	1623: sound1 <=  408569;
	1624: sound1 <=  376190;
	1625: sound1 <=  320038;
	1626: sound1 <=  230835;
	1627: sound1 <=  108215;
	1628: sound1 <=  2686;
	1629: sound1 <=  -58655;
	1630: sound1 <=  -118927;
	1631: sound1 <=  -154999;
	1632: sound1 <=  -149384;
	1633: sound1 <=  -170807;
	1634: sound1 <=  -200439;
	1635: sound1 <=  -233917;
	1636: sound1 <=  -257965;
	1637: sound1 <=  -286407;
	1638: sound1 <=  -323517;
	1639: sound1 <=  -326385;
	1640: sound1 <=  -323822;
	1641: sound1 <=  -311279;
	1642: sound1 <=  -312866;
	1643: sound1 <=  -258850;
	1644: sound1 <=  -197998;
	1645: sound1 <=  -193573;
	1646: sound1 <=  -173645;
	1647: sound1 <=  -148773;
	1648: sound1 <=  -137238;
	1649: sound1 <=  -123016;
	1650: sound1 <=  -102020;
	1651: sound1 <=  -80841;
	1652: sound1 <=  -29480;
	1653: sound1 <=  51270;
	1654: sound1 <=  116333;
	1655: sound1 <=  183105;
	1656: sound1 <=  246582;
	1657: sound1 <=  337982;
	1658: sound1 <=  420746;
	1659: sound1 <=  467926;
	1660: sound1 <=  505524;
	1661: sound1 <=  519501;
	1662: sound1 <=  517212;
	1663: sound1 <=  501404;
	1664: sound1 <=  451996;
	1665: sound1 <=  411072;
	1666: sound1 <=  402252;
	1667: sound1 <=  399231;
	1668: sound1 <=  389862;
	1669: sound1 <=  364044;
	1670: sound1 <=  329315;
	1671: sound1 <=  305084;
	1672: sound1 <=  288513;
	1673: sound1 <=  256042;
	1674: sound1 <=  235992;
	1675: sound1 <=  243500;
	1676: sound1 <=  232178;
	1677: sound1 <=  207581;
	1678: sound1 <=  220245;
	1679: sound1 <=  255951;
	1680: sound1 <=  274567;
	1681: sound1 <=  273438;
	1682: sound1 <=  269348;
	1683: sound1 <=  251801;
	1684: sound1 <=  214417;
	1685: sound1 <=  150330;
	1686: sound1 <=  33478;
	1687: sound1 <=  -94086;
	1688: sound1 <=  -217896;
	1689: sound1 <=  -329742;
	1690: sound1 <=  -398438;
	1691: sound1 <=  -429108;
	1692: sound1 <=  -408142;
	1693: sound1 <=  -377594;
	1694: sound1 <=  -354706;
	1695: sound1 <=  -308563;
	1696: sound1 <=  -286957;
	1697: sound1 <=  -289948;
	1698: sound1 <=  -315582;
	1699: sound1 <=  -318787;
	1700: sound1 <=  -332397;
	1701: sound1 <=  -388519;
	1702: sound1 <=  -402771;
	1703: sound1 <=  -395233;
	1704: sound1 <=  -386505;
	1705: sound1 <=  -386566;
	1706: sound1 <=  -390320;
	1707: sound1 <=  -373779;
	1708: sound1 <=  -351593;
	1709: sound1 <=  -341431;
	1710: sound1 <=  -307739;
	1711: sound1 <=  -231171;
	1712: sound1 <=  -169708;
	1713: sound1 <=  -105560;
	1714: sound1 <=  -47424;
	1715: sound1 <=  38971;
	1716: sound1 <=  114410;
	1717: sound1 <=  147064;
	1718: sound1 <=  171692;
	1719: sound1 <=  170654;
	1720: sound1 <=  139191;
	1721: sound1 <=  86121;
	1722: sound1 <=  33295;
	1723: sound1 <=  15198;
	1724: sound1 <=  -6744;
	1725: sound1 <=  -34271;
	1726: sound1 <=  -62134;
	1727: sound1 <=  -73334;
	1728: sound1 <=  -92560;
	1729: sound1 <=  -89752;
	1730: sound1 <=  -66986;
	1731: sound1 <=  -67657;
	1732: sound1 <=  -83130;
	1733: sound1 <=  -99274;
	1734: sound1 <=  -126160;
	1735: sound1 <=  -137329;
	1736: sound1 <=  -149780;
	1737: sound1 <=  -182007;
	1738: sound1 <=  -151947;
	1739: sound1 <=  -103760;
	1740: sound1 <=  -70740;
	1741: sound1 <=  -4700;
	1742: sound1 <=  76660;
	1743: sound1 <=  125763;
	1744: sound1 <=  137085;
	1745: sound1 <=  126099;
	1746: sound1 <=  146332;
	1747: sound1 <=  196777;
	1748: sound1 <=  235687;
	1749: sound1 <=  249573;
	1750: sound1 <=  304718;
	1751: sound1 <=  203430;
	1752: sound1 <=  -16357;
	1753: sound1 <=  2869;
	1754: sound1 <=  -8972;
	1755: sound1 <=  -4517;
	1756: sound1 <=  -6683;
	1757: sound1 <=  10681;
	1758: sound1 <=  36407;
	1759: sound1 <=  43854;
	1760: sound1 <=  66284;
	1761: sound1 <=  142853;
	1762: sound1 <=  196503;
	1763: sound1 <=  223480;
	1764: sound1 <=  276581;
	1765: sound1 <=  300934;
	1766: sound1 <=  341034;
	1767: sound1 <=  396790;
	1768: sound1 <=  464355;
	1769: sound1 <=  466003;
	1770: sound1 <=  441772;
	1771: sound1 <=  446655;
	1772: sound1 <=  441498;
	1773: sound1 <=  439484;
	1774: sound1 <=  450195;
	1775: sound1 <=  461670;
	1776: sound1 <=  456940;
	1777: sound1 <=  440887;
	1778: sound1 <=  424133;
	1779: sound1 <=  419342;
	1780: sound1 <=  412415;
	1781: sound1 <=  389954;
	1782: sound1 <=  356140;
	1783: sound1 <=  311890;
	1784: sound1 <=  239594;
	1785: sound1 <=  144928;
	1786: sound1 <=  67474;
	1787: sound1 <=  19531;
	1788: sound1 <=  -69397;
	1789: sound1 <=  -184662;
	1790: sound1 <=  -267670;
	1791: sound1 <=  -289856;
	1792: sound1 <=  -298981;
	1793: sound1 <=  -309082;
	1794: sound1 <=  -321411;
	1795: sound1 <=  -346527;
	1796: sound1 <=  -341309;
	1797: sound1 <=  -313751;
	1798: sound1 <=  -295898;
	1799: sound1 <=  -271149;
	1800: sound1 <=  -256958;
	1801: sound1 <=  -238678;
	1802: sound1 <=  -200317;
	1803: sound1 <=  -131531;
	1804: sound1 <=  -125824;
	1805: sound1 <=  -120270;
	1806: sound1 <=  -128082;
	1807: sound1 <=  -149109;
	1808: sound1 <=  -170410;
	1809: sound1 <=  -195709;
	1810: sound1 <=  -202423;
	1811: sound1 <=  -216187;
	1812: sound1 <=  -235962;
	1813: sound1 <=  -250153;
	1814: sound1 <=  -262543;
	1815: sound1 <=  -269379;
	1816: sound1 <=  -221863;
	1817: sound1 <=  -160187;
	1818: sound1 <=  -109863;
	1819: sound1 <=  -12146;
	1820: sound1 <=  45013;
	1821: sound1 <=  102753;
	1822: sound1 <=  163055;
	1823: sound1 <=  239044;
	1824: sound1 <=  289551;
	1825: sound1 <=  324219;
	1826: sound1 <=  363068;
	1827: sound1 <=  348297;
	1828: sound1 <=  358643;
	1829: sound1 <=  283386;
	1830: sound1 <=  57922;
	1831: sound1 <=  22705;
	1832: sound1 <=  -55603;
	1833: sound1 <=  -150146;
	1834: sound1 <=  -198456;
	1835: sound1 <=  -216400;
	1836: sound1 <=  -202698;
	1837: sound1 <=  -182922;
	1838: sound1 <=  -175354;
	1839: sound1 <=  -169983;
	1840: sound1 <=  -179779;
	1841: sound1 <=  -169830;
	1842: sound1 <=  -163177;
	1843: sound1 <=  -154724;
	1844: sound1 <=  -118561;
	1845: sound1 <=  -81879;
	1846: sound1 <=  -30060;
	1847: sound1 <=  48798;
	1848: sound1 <=  134979;
	1849: sound1 <=  184235;
	1850: sound1 <=  229584;
	1851: sound1 <=  305969;
	1852: sound1 <=  380524;
	1853: sound1 <=  441895;
	1854: sound1 <=  495422;
	1855: sound1 <=  552917;
	1856: sound1 <=  589935;
	1857: sound1 <=  587982;
	1858: sound1 <=  571564;
	1859: sound1 <=  509338;
	1860: sound1 <=  461761;
	1861: sound1 <=  420624;
	1862: sound1 <=  384766;
	1863: sound1 <=  321350;
	1864: sound1 <=  261505;
	1865: sound1 <=  193787;
	1866: sound1 <=  136688;
	1867: sound1 <=  82123;
	1868: sound1 <=  77209;
	1869: sound1 <=  46112;
	1870: sound1 <=  27588;
	1871: sound1 <=  -177094;
	1872: sound1 <=  -276947;
	1873: sound1 <=  -262299;
	1874: sound1 <=  -304626;
	1875: sound1 <=  -281647;
	1876: sound1 <=  -415741;
	1877: sound1 <=  -479645;
	1878: sound1 <=  -455597;
	1879: sound1 <=  -466095;
	1880: sound1 <=  -403381;
	1881: sound1 <=  -293762;
	1882: sound1 <=  -249939;
	1883: sound1 <=  -304382;
	1884: sound1 <=  -263275;
	1885: sound1 <=  -256165;
	1886: sound1 <=  -230042;
	1887: sound1 <=  -208038;
	1888: sound1 <=  -201172;
	1889: sound1 <=  -185730;
	1890: sound1 <=  -167999;
	1891: sound1 <=  -155609;
	1892: sound1 <=  -141724;
	1893: sound1 <=  -121399;
	1894: sound1 <=  -88318;
	1895: sound1 <=  -52307;
	1896: sound1 <=  -1312;
	1897: sound1 <=  50446;
	1898: sound1 <=  71564;
	1899: sound1 <=  74707;
	1900: sound1 <=  74402;
	1901: sound1 <=  82123;
	1902: sound1 <=  80017;
	1903: sound1 <=  59753;
	1904: sound1 <=  31189;
	1905: sound1 <=  33295;
	1906: sound1 <=  48218;
	1907: sound1 <=  62347;
	1908: sound1 <=  92560;
	1909: sound1 <=  125946;
	1910: sound1 <=  124084;
	1911: sound1 <=  124451;
	1912: sound1 <=  120605;
	1913: sound1 <=  119446;
	1914: sound1 <=  151764;
	1915: sound1 <=  222839;
	1916: sound1 <=  197571;
	1917: sound1 <=  -31555;
	1918: sound1 <=  -64056;
	1919: sound1 <=  -39581;
	1920: sound1 <=  -45898;
	1921: sound1 <=  -64026;
	1922: sound1 <=  -90698;
	1923: sound1 <=  -67169;
	1924: sound1 <=  -88074;
	1925: sound1 <=  -108856;
	1926: sound1 <=  -116760;
	1927: sound1 <=  -138641;
	1928: sound1 <=  -125580;
	1929: sound1 <=  -113098;
	1930: sound1 <=  -58350;
	1931: sound1 <=  -61;
	1932: sound1 <=  55389;
	1933: sound1 <=  156433;
	1934: sound1 <=  263824;
	1935: sound1 <=  350586;
	1936: sound1 <=  409119;
	1937: sound1 <=  472198;
	1938: sound1 <=  549988;
	1939: sound1 <=  637848;
	1940: sound1 <=  670471;
	1941: sound1 <=  661926;
	1942: sound1 <=  646698;
	1943: sound1 <=  598206;
	1944: sound1 <=  552216;
	1945: sound1 <=  524597;
	1946: sound1 <=  492950;
	1947: sound1 <=  450836;
	1948: sound1 <=  399811;
	1949: sound1 <=  326813;
	1950: sound1 <=  241241;
	1951: sound1 <=  184387;
	1952: sound1 <=  142487;
	1953: sound1 <=  102814;
	1954: sound1 <=  80841;
	1955: sound1 <=  62469;
	1956: sound1 <=  56580;
	1957: sound1 <=  43549;
	1958: sound1 <=  20569;
	1959: sound1 <=  4852;
	1960: sound1 <=  -26886;
	1961: sound1 <=  -52521;
	1962: sound1 <=  -52185;
	1963: sound1 <=  -33691;
	1964: sound1 <=  -15900;
	1965: sound1 <=  -28534;
	1966: sound1 <=  -70435;
	1967: sound1 <=  -130585;
	1968: sound1 <=  -114685;
	1969: sound1 <=  -67535;
	1970: sound1 <=  -47852;
	1971: sound1 <=  -49957;
	1972: sound1 <=  -79620;
	1973: sound1 <=  -103241;
	1974: sound1 <=  -118713;
	1975: sound1 <=  -141876;
	1976: sound1 <=  -163116;
	1977: sound1 <=  -194794;
	1978: sound1 <=  -217194;
	1979: sound1 <=  -228271;
	1980: sound1 <=  -231293;
	1981: sound1 <=  -257141;
	1982: sound1 <=  -268127;
	1983: sound1 <=  -283386;
	1984: sound1 <=  -311554;
	1985: sound1 <=  -301483;
	1986: sound1 <=  -290833;
	1987: sound1 <=  -287415;
	1988: sound1 <=  -283875;
	1989: sound1 <=  -290192;
	1990: sound1 <=  -281799;
	1991: sound1 <=  -248810;
	1992: sound1 <=  -224792;
	1993: sound1 <=  -229492;
	1994: sound1 <=  -186432;
	1995: sound1 <=  -162994;
	1996: sound1 <=  -137482;
	1997: sound1 <=  -116821;
	1998: sound1 <=  -85449;
	1999: sound1 <=  -36896;
	2000: sound1 <=  -12512;
	2001: sound1 <=  32990;
	2002: sound1 <=  72266;
	2003: sound1 <=  65460;
	2004: sound1 <=  94666;
	2005: sound1 <=  157471;
	2006: sound1 <=  189117;
	2007: sound1 <=  204376;
	2008: sound1 <=  205444;
	2009: sound1 <=  216278;
	2010: sound1 <=  204926;
	2011: sound1 <=  144531;
	2012: sound1 <=  -67780;
	2013: sound1 <=  -123016;
	2014: sound1 <=  -102356;
	2015: sound1 <=  -103821;
	2016: sound1 <=  -90668;
	2017: sound1 <=  -79193;
	2018: sound1 <=  -66193;
	2019: sound1 <=  -57373;
	2020: sound1 <=  -60455;
	2021: sound1 <=  -89081;
	2022: sound1 <=  -98419;
	2023: sound1 <=  -108154;
	2024: sound1 <=  -116730;
	2025: sound1 <=  -100891;
	2026: sound1 <=  -83649;
	2027: sound1 <=  -80933;
	2028: sound1 <=  -45105;
	2029: sound1 <=  -2899;
	2030: sound1 <=  63263;
	2031: sound1 <=  142761;
	2032: sound1 <=  219452;
	2033: sound1 <=  286591;
	2034: sound1 <=  328369;
	2035: sound1 <=  359283;
	2036: sound1 <=  352509;
	2037: sound1 <=  357483;
	2038: sound1 <=  398071;
	2039: sound1 <=  432678;
	2040: sound1 <=  449219;
	2041: sound1 <=  435394;
	2042: sound1 <=  441376;
	2043: sound1 <=  447174;
	2044: sound1 <=  451965;
	2045: sound1 <=  428986;
	2046: sound1 <=  401550;
	2047: sound1 <=  367340;
	2048: sound1 <=  323639;
	2049: sound1 <=  293884;
	2050: sound1 <=  241089;
	2051: sound1 <=  169281;
	2052: sound1 <=  120514;
	2053: sound1 <=  48279;
	2054: sound1 <=  -39703;
	2055: sound1 <=  -131836;
	2056: sound1 <=  -225037;
	2057: sound1 <=  -238922;
	2058: sound1 <=  -248749;
	2059: sound1 <=  -284241;
	2060: sound1 <=  -312500;
	2061: sound1 <=  -335266;
	2062: sound1 <=  -315674;
	2063: sound1 <=  -295471;
	2064: sound1 <=  -261749;
	2065: sound1 <=  -268890;
	2066: sound1 <=  -275726;
	2067: sound1 <=  -268036;
	2068: sound1 <=  -246521;
	2069: sound1 <=  -210358;
	2070: sound1 <=  -202057;
	2071: sound1 <=  -212494;
	2072: sound1 <=  -200226;
	2073: sound1 <=  -152100;
	2074: sound1 <=  -76691;
	2075: sound1 <=  2136;
	2076: sound1 <=  109589;
	2077: sound1 <=  180298;
	2078: sound1 <=  270142;
	2079: sound1 <=  346588;
	2080: sound1 <=  405762;
	2081: sound1 <=  453552;
	2082: sound1 <=  468842;
	2083: sound1 <=  440277;
	2084: sound1 <=  391174;
	2085: sound1 <=  375824;
	2086: sound1 <=  376129;
	2087: sound1 <=  361450;
	2088: sound1 <=  345001;
	2089: sound1 <=  341736;
	2090: sound1 <=  311829;
	2091: sound1 <=  283447;
	2092: sound1 <=  177612;
	2093: sound1 <=  120728;
	2094: sound1 <=  178619;
	2095: sound1 <=  87402;
	2096: sound1 <=  -32318;
	2097: sound1 <=  -45288;
	2098: sound1 <=  -108826;
	2099: sound1 <=  -143738;
	2100: sound1 <=  -186859;
	2101: sound1 <=  -198792;
	2102: sound1 <=  -133636;
	2103: sound1 <=  -192352;
	2104: sound1 <=  -243164;
	2105: sound1 <=  -179169;
	2106: sound1 <=  -181122;
	2107: sound1 <=  -197906;
	2108: sound1 <=  -188721;
	2109: sound1 <=  -201019;
	2110: sound1 <=  -186829;
	2111: sound1 <=  -168732;
	2112: sound1 <=  -206177;
	2113: sound1 <=  -237091;
	2114: sound1 <=  -197174;
	2115: sound1 <=  -103424;
	2116: sound1 <=  -81757;
	2117: sound1 <=  -107422;
	2118: sound1 <=  22461;
	2119: sound1 <=  -54321;
	2120: sound1 <=  27557;
	2121: sound1 <=  93536;
	2122: sound1 <=  20660;
	2123: sound1 <=  98450;
	2124: sound1 <=  133514;
	2125: sound1 <=  -31525;
	2126: sound1 <=  -76385;
	2127: sound1 <=  -39825;
	2128: sound1 <=  -18738;
	2129: sound1 <=  -8179;
	2130: sound1 <=  -138519;
	2131: sound1 <=  -61096;
	2132: sound1 <=  -3693;
	2133: sound1 <=  -26459;
	2134: sound1 <=  -21912;
	2135: sound1 <=  -169342;
	2136: sound1 <=  -143585;
	2137: sound1 <=  -134949;
	2138: sound1 <=  -59723;
	2139: sound1 <=  -118195;
	2140: sound1 <=  -69824;
	2141: sound1 <=  -92560;
	2142: sound1 <=  -60638;
	2143: sound1 <=  -78735;
	2144: sound1 <=  -44739;
	2145: sound1 <=  -66742;
	2146: sound1 <=  -38666;
	2147: sound1 <=  61951;
	2148: sound1 <=  125916;
	2149: sound1 <=  -11200;
	2150: sound1 <=  -133514;
	2151: sound1 <=  -71533;
	2152: sound1 <=  -41656;
	2153: sound1 <=  28778;
	2154: sound1 <=  98236;
	2155: sound1 <=  127502;
	2156: sound1 <=  169403;
	2157: sound1 <=  183838;
	2158: sound1 <=  193665;
	2159: sound1 <=  51422;
	2160: sound1 <=  -3998;
	2161: sound1 <=  21942;
	2162: sound1 <=  68878;
	2163: sound1 <=  144897;
	2164: sound1 <=  236877;
	2165: sound1 <=  229187;
	2166: sound1 <=  161407;
	2167: sound1 <=  226563;
	2168: sound1 <=  277130;
	2169: sound1 <=  246552;
	2170: sound1 <=  250641;
	2171: sound1 <=  306091;
	2172: sound1 <=  337982;
	2173: sound1 <=  256256;
	2174: sound1 <=  157837;
	2175: sound1 <=  153351;
	2176: sound1 <=  120880;
	2177: sound1 <=  150848;
	2178: sound1 <=  131836;
	2179: sound1 <=  158356;
	2180: sound1 <=  215851;
	2181: sound1 <=  272003;
	2182: sound1 <=  308197;
	2183: sound1 <=  343933;
	2184: sound1 <=  239014;
	2185: sound1 <=  250580;
	2186: sound1 <=  278442;
	2187: sound1 <=  278168;
	2188: sound1 <=  281677;
	2189: sound1 <=  234070;
	2190: sound1 <=  203430;
	2191: sound1 <=  3418;
	2192: sound1 <=  -112762;
	2193: sound1 <=  -101501;
	2194: sound1 <=  -104065;
	2195: sound1 <=  -109436;
	2196: sound1 <=  -69824;
	2197: sound1 <=  -14069;
	2198: sound1 <=  55054;
	2199: sound1 <=  12115;
	2200: sound1 <=  -173828;
	2201: sound1 <=  -113617;
	2202: sound1 <=  -121002;
	2203: sound1 <=  -139801;
	2204: sound1 <=  -177917;
	2205: sound1 <=  -160339;
	2206: sound1 <=  -134918;
	2207: sound1 <=  -113739;
	2208: sound1 <=  -68268;
	2209: sound1 <=  -21240;
	2210: sound1 <=  50934;
	2211: sound1 <=  130524;
	2212: sound1 <=  170258;
	2213: sound1 <=  183502;
	2214: sound1 <=  185577;
	2215: sound1 <=  196075;
	2216: sound1 <=  159363;
	2217: sound1 <=  139832;
	2218: sound1 <=  140717;
	2219: sound1 <=  101318;
	2220: sound1 <=  83191;
	2221: sound1 <=  46753;
	2222: sound1 <=  32623;
	2223: sound1 <=  -171814;
	2224: sound1 <=  -370026;
	2225: sound1 <=  -339386;
	2226: sound1 <=  -320740;
	2227: sound1 <=  -295746;
	2228: sound1 <=  -279633;
	2229: sound1 <=  -239471;
	2230: sound1 <=  -202301;
	2231: sound1 <=  -187988;
	2232: sound1 <=  -166595;
	2233: sound1 <=  -120422;
	2234: sound1 <=  -64545;
	2235: sound1 <=  25391;
	2236: sound1 <=  143066;
	2237: sound1 <=  178040;
	2238: sound1 <=  195801;
	2239: sound1 <=  53558;
	2240: sound1 <=  15289;
	2241: sound1 <=  62317;
	2242: sound1 <=  99335;
	2243: sound1 <=  186523;
	2244: sound1 <=  212860;
	2245: sound1 <=  213837;
	2246: sound1 <=  197784;
	2247: sound1 <=  192780;
	2248: sound1 <=  153351;
	2249: sound1 <=  99548;
	2250: sound1 <=  40009;
	2251: sound1 <=  7141;
	2252: sound1 <=  -6317;
	2253: sound1 <=  -31097;
	2254: sound1 <=  -18219;
	2255: sound1 <=  12726;
	2256: sound1 <=  9033;
	2257: sound1 <=  14862;
	2258: sound1 <=  23010;
	2259: sound1 <=  62378;
	2260: sound1 <=  46021;
	2261: sound1 <=  4242;
	2262: sound1 <=  -458;
	2263: sound1 <=  -35980;
	2264: sound1 <=  -65674;
	2265: sound1 <=  -92438;
	2266: sound1 <=  -106354;
	2267: sound1 <=  -113953;
	2268: sound1 <=  -91766;
	2269: sound1 <=  -70740;
	2270: sound1 <=  -78094;
	2271: sound1 <=  -92590;
	2272: sound1 <=  -110199;
	2273: sound1 <=  -150085;
	2274: sound1 <=  -147888;
	2275: sound1 <=  -90179;
	2276: sound1 <=  -73944;
	2277: sound1 <=  -90149;
	2278: sound1 <=  -118500;
	2279: sound1 <=  -124359;
	2280: sound1 <=  -101929;
	2281: sound1 <=  -84900;
	2282: sound1 <=  -105133;
	2283: sound1 <=  -115326;
	2284: sound1 <=  -103882;
	2285: sound1 <=  -75043;
	2286: sound1 <=  -47821;
	2287: sound1 <=  -23712;
	2288: sound1 <=  16693;
	2289: sound1 <=  104401;
	2290: sound1 <=  198975;
	2291: sound1 <=  292114;
	2292: sound1 <=  333679;
	2293: sound1 <=  355255;
	2294: sound1 <=  364502;
	2295: sound1 <=  373779;
	2296: sound1 <=  374786;
	2297: sound1 <=  372650;
	2298: sound1 <=  377441;
	2299: sound1 <=  379242;
	2300: sound1 <=  338745;
	2301: sound1 <=  301666;
	2302: sound1 <=  293701;
	2303: sound1 <=  303467;
	2304: sound1 <=  318237;
	2305: sound1 <=  299347;
	2306: sound1 <=  275208;
	2307: sound1 <=  271210;
	2308: sound1 <=  269531;
	2309: sound1 <=  243988;
	2310: sound1 <=  210693;
	2311: sound1 <=  165253;
	2312: sound1 <=  134705;
	2313: sound1 <=  141052;
	2314: sound1 <=  123077;
	2315: sound1 <=  105804;
	2316: sound1 <=  92194;
	2317: sound1 <=  71747;
	2318: sound1 <=  24200;
	2319: sound1 <=  -46814;
	2320: sound1 <=  -73364;
	2321: sound1 <=  -68542;
	2322: sound1 <=  -56000;
	2323: sound1 <=  -37750;
	2324: sound1 <=  5005;
	2325: sound1 <=  49286;
	2326: sound1 <=  82886;
	2327: sound1 <=  73395;
	2328: sound1 <=  59448;
	2329: sound1 <=  56580;
	2330: sound1 <=  44312;
	2331: sound1 <=  38849;
	2332: sound1 <=  16052;
	2333: sound1 <=  -21515;
	2334: sound1 <=  -54474;
	2335: sound1 <=  -40955;
	2336: sound1 <=  -116577;
	2337: sound1 <=  -333405;
	2338: sound1 <=  -327271;
	2339: sound1 <=  -344543;
	2340: sound1 <=  -373047;
	2341: sound1 <=  -372162;
	2342: sound1 <=  -357086;
	2343: sound1 <=  -340851;
	2344: sound1 <=  -316498;
	2345: sound1 <=  -294678;
	2346: sound1 <=  -273834;
	2347: sound1 <=  -244781;
	2348: sound1 <=  -221161;
	2349: sound1 <=  -217529;
	2350: sound1 <=  -188385;
	2351: sound1 <=  -151703;
	2352: sound1 <=  -133942;
	2353: sound1 <=  -188660;
	2354: sound1 <=  -224243;
	2355: sound1 <=  -243347;
	2356: sound1 <=  -251709;
	2357: sound1 <=  -239288;
	2358: sound1 <=  -263855;
	2359: sound1 <=  -274200;
	2360: sound1 <=  -249023;
	2361: sound1 <=  -247772;
	2362: sound1 <=  -238434;
	2363: sound1 <=  -234741;
	2364: sound1 <=  -217865;
	2365: sound1 <=  -178467;
	2366: sound1 <=  -202698;
	2367: sound1 <=  -201721;
	2368: sound1 <=  -125092;
	2369: sound1 <=  -30029;
	2370: sound1 <=  38574;
	2371: sound1 <=  86212;
	2372: sound1 <=  115814;
	2373: sound1 <=  143127;
	2374: sound1 <=  164215;
	2375: sound1 <=  195068;
	2376: sound1 <=  202148;
	2377: sound1 <=  192352;
	2378: sound1 <=  212830;
	2379: sound1 <=  249603;
	2380: sound1 <=  273102;
	2381: sound1 <=  278809;
	2382: sound1 <=  313751;
	2383: sound1 <=  329407;
	2384: sound1 <=  334290;
	2385: sound1 <=  302246;
	2386: sound1 <=  278625;
	2387: sound1 <=  269653;
	2388: sound1 <=  295410;
	2389: sound1 <=  308411;
	2390: sound1 <=  282257;
	2391: sound1 <=  258972;
	2392: sound1 <=  230835;
	2393: sound1 <=  224182;
	2394: sound1 <=  221771;
	2395: sound1 <=  219543;
	2396: sound1 <=  205078;
	2397: sound1 <=  205688;
	2398: sound1 <=  211121;
	2399: sound1 <=  188324;
	2400: sound1 <=  142578;
	2401: sound1 <=  112518;
	2402: sound1 <=  118378;
	2403: sound1 <=  133240;
	2404: sound1 <=  130951;
	2405: sound1 <=  140076;
	2406: sound1 <=  159668;
	2407: sound1 <=  192108;
	2408: sound1 <=  235809;
	2409: sound1 <=  278046;
	2410: sound1 <=  276917;
	2411: sound1 <=  268280;
	2412: sound1 <=  90454;
	2413: sound1 <=  44464;
	2414: sound1 <=  49438;
	2415: sound1 <=  9369;
	2416: sound1 <=  -36194;
	2417: sound1 <=  -78735;
	2418: sound1 <=  -57922;
	2419: sound1 <=  -75165;
	2420: sound1 <=  -68268;
	2421: sound1 <=  -26550;
	2422: sound1 <=  -27039;
	2423: sound1 <=  -181915;
	2424: sound1 <=  -163666;
	2425: sound1 <=  -140228;
	2426: sound1 <=  -151550;
	2427: sound1 <=  -95093;
	2428: sound1 <=  -16846;
	2429: sound1 <=  27435;
	2430: sound1 <=  75409;
	2431: sound1 <=  98267;
	2432: sound1 <=  116638;
	2433: sound1 <=  -37964;
	2434: sound1 <=  -184540;
	2435: sound1 <=  -185974;
	2436: sound1 <=  -186188;
	2437: sound1 <=  -179535;
	2438: sound1 <=  -158905;
	2439: sound1 <=  -134766;
	2440: sound1 <=  -87067;
	2441: sound1 <=  -58014;
	2442: sound1 <=  -35095;
	2443: sound1 <=  31311;
	2444: sound1 <=  120178;
	2445: sound1 <=  196960;
	2446: sound1 <=  140381;
	2447: sound1 <=  2533;
	2448: sound1 <=  19440;
	2449: sound1 <=  -12054;
	2450: sound1 <=  -11108;
	2451: sound1 <=  23224;
	2452: sound1 <=  48157;
	2453: sound1 <=  75897;
	2454: sound1 <=  96985;
	2455: sound1 <=  109131;
	2456: sound1 <=  147858;
	2457: sound1 <=  161530;
	2458: sound1 <=  138275;
	2459: sound1 <=  115326;
	2460: sound1 <=  101868;
	2461: sound1 <=  97046;
	2462: sound1 <=  121490;
	2463: sound1 <=  163727;
	2464: sound1 <=  197327;
	2465: sound1 <=  -153;
	2466: sound1 <=  -56488;
	2467: sound1 <=  -41809;
	2468: sound1 <=  -21637;
	2469: sound1 <=  -6775;
	2470: sound1 <=  9277;
	2471: sound1 <=  34851;
	2472: sound1 <=  12848;
	2473: sound1 <=  -13092;
	2474: sound1 <=  13794;
	2475: sound1 <=  84839;
	2476: sound1 <=  85663;
	2477: sound1 <=  108795;
	2478: sound1 <=  132538;
	2479: sound1 <=  191711;
	2480: sound1 <=  111816;
	2481: sound1 <=  -32990;
	2482: sound1 <=  -19806;
	2483: sound1 <=  -64087;
	2484: sound1 <=  -69275;
	2485: sound1 <=  -21149;
	2486: sound1 <=  36255;
	2487: sound1 <=  83527;
	2488: sound1 <=  142059;
	2489: sound1 <=  198029;
	2490: sound1 <=  219940;
	2491: sound1 <=  209015;
	2492: sound1 <=  179626;
	2493: sound1 <=  174255;
	2494: sound1 <=  -9644;
	2495: sound1 <=  -159882;
	2496: sound1 <=  -172607;
	2497: sound1 <=  -225189;
	2498: sound1 <=  -254486;
	2499: sound1 <=  -280640;
	2500: sound1 <=  -283173;
	2501: sound1 <=  -268311;
	2502: sound1 <=  -229065;
	2503: sound1 <=  -192688;
	2504: sound1 <=  -176178;
	2505: sound1 <=  -182190;
	2506: sound1 <=  -197540;
	2507: sound1 <=  -178925;
	2508: sound1 <=  -126312;
	2509: sound1 <=  -60059;
	2510: sound1 <=  4364;
	2511: sound1 <=  56641;
	2512: sound1 <=  50446;
	2513: sound1 <=  67963;
	2514: sound1 <=  130371;
	2515: sound1 <=  191132;
	2516: sound1 <=  295776;
	2517: sound1 <=  353088;
	2518: sound1 <=  349640;
	2519: sound1 <=  355255;
	2520: sound1 <=  390106;
	2521: sound1 <=  415497;
	2522: sound1 <=  427032;
	2523: sound1 <=  392487;
	2524: sound1 <=  348114;
	2525: sound1 <=  333435;
	2526: sound1 <=  342468;
	2527: sound1 <=  356262;
	2528: sound1 <=  369934;
	2529: sound1 <=  357208;
	2530: sound1 <=  311646;
	2531: sound1 <=  241516;
	2532: sound1 <=  204926;
	2533: sound1 <=  61554;
	2534: sound1 <=  -203003;
	2535: sound1 <=  -232239;
	2536: sound1 <=  -284332;
	2537: sound1 <=  -295441;
	2538: sound1 <=  -291901;
	2539: sound1 <=  -308136;
	2540: sound1 <=  -278351;
	2541: sound1 <=  -249359;
	2542: sound1 <=  -212250;
	2543: sound1 <=  -201935;
	2544: sound1 <=  -188446;
	2545: sound1 <=  -106537;
	2546: sound1 <=  -42450;
	2547: sound1 <=  -15961;
	2548: sound1 <=  -53101;
	2549: sound1 <=  -135315;
	2550: sound1 <=  -124725;
	2551: sound1 <=  -119019;
	2552: sound1 <=  -99548;
	2553: sound1 <=  -99335;
	2554: sound1 <=  -121643;
	2555: sound1 <=  -148193;
	2556: sound1 <=  -175354;
	2557: sound1 <=  -195526;
	2558: sound1 <=  -159698;
	2559: sound1 <=  -106293;
	2560: sound1 <=  -24719;
	2561: sound1 <=  29449;
	2562: sound1 <=  57831;
	2563: sound1 <=  83282;
	2564: sound1 <=  126984;
	2565: sound1 <=  139252;
	2566: sound1 <=  165039;
	2567: sound1 <=  184082;
	2568: sound1 <=  193298;
	2569: sound1 <=  214996;
	2570: sound1 <=  240021;
	2571: sound1 <=  154480;
	2572: sound1 <=  94635;
	2573: sound1 <=  143311;
	2574: sound1 <=  171875;
	2575: sound1 <=  181610;
	2576: sound1 <=  165619;
	2577: sound1 <=  160858;
	2578: sound1 <=  120972;
	2579: sound1 <=  99365;
	2580: sound1 <=  84808;
	2581: sound1 <=  -136963;
	2582: sound1 <=  -194214;
	2583: sound1 <=  -233093;
	2584: sound1 <=  -247833;
	2585: sound1 <=  -194672;
	2586: sound1 <=  -141785;
	2587: sound1 <=  -94391;
	2588: sound1 <=  -76355;
	2589: sound1 <=  -67719;
	2590: sound1 <=  -56671;
	2591: sound1 <=  -79559;
	2592: sound1 <=  -59998;
	2593: sound1 <=  -26306;
	2594: sound1 <=  -20752;
	2595: sound1 <=  -10254;
	2596: sound1 <=  54352;
	2597: sound1 <=  117737;
	2598: sound1 <=  194458;
	2599: sound1 <=  233795;
	2600: sound1 <=  258209;
	2601: sound1 <=  280121;
	2602: sound1 <=  271057;
	2603: sound1 <=  297119;
	2604: sound1 <=  311066;
	2605: sound1 <=  282318;
	2606: sound1 <=  193542;
	2607: sound1 <=  -67352;
	2608: sound1 <=  -166718;
	2609: sound1 <=  -215240;
	2610: sound1 <=  -214569;
	2611: sound1 <=  -219238;
	2612: sound1 <=  -247650;
	2613: sound1 <=  -260864;
	2614: sound1 <=  -256897;
	2615: sound1 <=  -268097;
	2616: sound1 <=  -249023;
	2617: sound1 <=  -231567;
	2618: sound1 <=  -232727;
	2619: sound1 <=  -186188;
	2620: sound1 <=  -150757;
	2621: sound1 <=  -117584;
	2622: sound1 <=  -92773;
	2623: sound1 <=  -28198;
	2624: sound1 <=  41260;
	2625: sound1 <=  66162;
	2626: sound1 <=  74188;
	2627: sound1 <=  98328;
	2628: sound1 <=  128265;
	2629: sound1 <=  184875;
	2630: sound1 <=  265228;
	2631: sound1 <=  282715;
	2632: sound1 <=  326782;
	2633: sound1 <=  373474;
	2634: sound1 <=  370789;
	2635: sound1 <=  395996;
	2636: sound1 <=  405396;
	2637: sound1 <=  396820;
	2638: sound1 <=  408997;
	2639: sound1 <=  397461;
	2640: sound1 <=  378632;
	2641: sound1 <=  367859;
	2642: sound1 <=  341400;
	2643: sound1 <=  326538;
	2644: sound1 <=  307220;
	2645: sound1 <=  310394;
	2646: sound1 <=  297119;
	2647: sound1 <=  278442;
	2648: sound1 <=  211548;
	2649: sound1 <=  157623;
	2650: sound1 <=  127228;
	2651: sound1 <=  108154;
	2652: sound1 <=  104950;
	2653: sound1 <=  100647;
	2654: sound1 <=  99304;
	2655: sound1 <=  91919;
	2656: sound1 <=  87372;
	2657: sound1 <=  27252;
	2658: sound1 <=  10773;
	2659: sound1 <=  6592;
	2660: sound1 <=  -21515;
	2661: sound1 <=  -52399;
	2662: sound1 <=  -79620;
	2663: sound1 <=  -109344;
	2664: sound1 <=  -149078;
	2665: sound1 <=  -157776;
	2666: sound1 <=  -170135;
	2667: sound1 <=  -154266;
	2668: sound1 <=  -133575;
	2669: sound1 <=  -149963;
	2670: sound1 <=  -162140;
	2671: sound1 <=  -187561;
	2672: sound1 <=  -227417;
	2673: sound1 <=  -229187;
	2674: sound1 <=  -248505;
	2675: sound1 <=  -300842;
	2676: sound1 <=  -307129;
	2677: sound1 <=  -298492;
	2678: sound1 <=  -299652;
	2679: sound1 <=  -296326;
	2680: sound1 <=  -312927;
	2681: sound1 <=  -313354;
	2682: sound1 <=  -307892;
	2683: sound1 <=  -317413;
	2684: sound1 <=  -282776;
	2685: sound1 <=  -250092;
	2686: sound1 <=  -223724;
	2687: sound1 <=  -200806;
	2688: sound1 <=  -211334;
	2689: sound1 <=  -171570;
	2690: sound1 <=  -140564;
	2691: sound1 <=  -97321;
	2692: sound1 <=  -55328;
	2693: sound1 <=  -40863;
	2694: sound1 <=  -17059;
	2695: sound1 <=  21271;
	2696: sound1 <=  20416;
	2697: sound1 <=  25391;
	2698: sound1 <=  32745;
	2699: sound1 <=  30029;
	2700: sound1 <=  3540;
	2701: sound1 <=  -43732;
	2702: sound1 <=  -32227;
	2703: sound1 <=  -8270;
	2704: sound1 <=  -9338;
	2705: sound1 <=  -11841;
	2706: sound1 <=  -45959;
	2707: sound1 <=  -52856;
	2708: sound1 <=  -48431;
	2709: sound1 <=  -57770;
	2710: sound1 <=  -30640;
	2711: sound1 <=  -9216;
	2712: sound1 <=  2594;
	2713: sound1 <=  61066;
	2714: sound1 <=  108551;
	2715: sound1 <=  146423;
	2716: sound1 <=  173492;
	2717: sound1 <=  177155;
	2718: sound1 <=  207123;
	2719: sound1 <=  230072;
	2720: sound1 <=  236877;
	2721: sound1 <=  231689;
	2722: sound1 <=  216339;
	2723: sound1 <=  260040;
	2724: sound1 <=  287018;
	2725: sound1 <=  271729;
	2726: sound1 <=  287903;
	2727: sound1 <=  323853;
	2728: sound1 <=  375854;
	2729: sound1 <=  399048;
	2730: sound1 <=  384125;
	2731: sound1 <=  374298;
	2732: sound1 <=  328918;
	2733: sound1 <=  288757;
	2734: sound1 <=  272919;
	2735: sound1 <=  231293;
	2736: sound1 <=  155273;
	2737: sound1 <=  135010;
	2738: sound1 <=  92255;
	2739: sound1 <=  60913;
	2740: sound1 <=  12451;
	2741: sound1 <=  -14282;
	2742: sound1 <=  -28931;
	2743: sound1 <=  -26245;
	2744: sound1 <=  -25635;
	2745: sound1 <=  -62775;
	2746: sound1 <=  -125000;
	2747: sound1 <=  -121613;
	2748: sound1 <=  -85236;
	2749: sound1 <=  -63507;
	2750: sound1 <=  -66345;
	2751: sound1 <=  -99121;
	2752: sound1 <=  -94177;
	2753: sound1 <=  -113556;
	2754: sound1 <=  -157837;
	2755: sound1 <=  -167358;
	2756: sound1 <=  -158997;
	2757: sound1 <=  -114868;
	2758: sound1 <=  -48645;
	2759: sound1 <=  -57037;
	2760: sound1 <=  -47058;
	2761: sound1 <=  34546;
	2762: sound1 <=  84778;
	2763: sound1 <=  147736;
	2764: sound1 <=  153564;
	2765: sound1 <=  142609;
	2766: sound1 <=  98267;
	2767: sound1 <=  75806;
	2768: sound1 <=  82977;
	2769: sound1 <=  88837;
	2770: sound1 <=  52643;
	2771: sound1 <=  34271;
	2772: sound1 <=  4669;
	2773: sound1 <=  -26154;
	2774: sound1 <=  -10590;
	2775: sound1 <=  -23346;
	2776: sound1 <=  1282;
	2777: sound1 <=  9766;
	2778: sound1 <=  -15503;
	2779: sound1 <=  -60486;
	2780: sound1 <=  -69183;
	2781: sound1 <=  -55145;
	2782: sound1 <=  -80719;
	2783: sound1 <=  -86212;
	2784: sound1 <=  -103394;
	2785: sound1 <=  -102264;
	2786: sound1 <=  -66498;
	2787: sound1 <=  -43762;
	2788: sound1 <=  -67505;
	2789: sound1 <=  -105225;
	2790: sound1 <=  -121826;
	2791: sound1 <=  -123596;
	2792: sound1 <=  -115417;
	2793: sound1 <=  -151550;
	2794: sound1 <=  -196899;
	2795: sound1 <=  -223206;
	2796: sound1 <=  -210022;
	2797: sound1 <=  -173553;
	2798: sound1 <=  -153839;
	2799: sound1 <=  -137482;
	2800: sound1 <=  -57922;
	2801: sound1 <=  31433;
	2802: sound1 <=  115540;
	2803: sound1 <=  171204;
	2804: sound1 <=  212250;
	2805: sound1 <=  269165;
	2806: sound1 <=  312927;
	2807: sound1 <=  377594;
	2808: sound1 <=  455231;
	2809: sound1 <=  493896;
	2810: sound1 <=  528320;
	2811: sound1 <=  591309;
	2812: sound1 <=  587341;
	2813: sound1 <=  541870;
	2814: sound1 <=  525726;
	2815: sound1 <=  510773;
	2816: sound1 <=  500641;
	2817: sound1 <=  500366;
	2818: sound1 <=  501434;
	2819: sound1 <=  498077;
	2820: sound1 <=  480072;
	2821: sound1 <=  437408;
	2822: sound1 <=  400299;
	2823: sound1 <=  397034;
	2824: sound1 <=  381744;
	2825: sound1 <=  349213;
	2826: sound1 <=  333221;
	2827: sound1 <=  315491;
	2828: sound1 <=  314545;
	2829: sound1 <=  288818;
	2830: sound1 <=  259430;
	2831: sound1 <=  229218;
	2832: sound1 <=  203979;
	2833: sound1 <=  205627;
	2834: sound1 <=  198090;
	2835: sound1 <=  146515;
	2836: sound1 <=  99030;
	2837: sound1 <=  55786;
	2838: sound1 <=  43121;
	2839: sound1 <=  44525;
	2840: sound1 <=  17426;
	2841: sound1 <=  9277;
	2842: sound1 <=  -10864;
	2843: sound1 <=  11993;
	2844: sound1 <=  49896;
	2845: sound1 <=  53284;
	2846: sound1 <=  18097;
	2847: sound1 <=  -33417;
	2848: sound1 <=  -70862;
	2849: sound1 <=  -49927;
	2850: sound1 <=  -39917;
	2851: sound1 <=  -95306;
	2852: sound1 <=  -136353;
	2853: sound1 <=  -196594;
	2854: sound1 <=  -218414;
	2855: sound1 <=  -228180;
	2856: sound1 <=  -267975;
	2857: sound1 <=  -301025;
	2858: sound1 <=  -329071;
	2859: sound1 <=  -332855;
	2860: sound1 <=  -339447;
	2861: sound1 <=  -340424;
	2862: sound1 <=  -320923;
	2863: sound1 <=  -316254;
	2864: sound1 <=  -409851;
	2865: sound1 <=  -418884;
	2866: sound1 <=  -430389;
	2867: sound1 <=  -431335;
	2868: sound1 <=  -419830;
	2869: sound1 <=  -436646;
	2870: sound1 <=  -441956;
	2871: sound1 <=  -466736;
	2872: sound1 <=  -478180;
	2873: sound1 <=  -472321;
	2874: sound1 <=  -444702;
	2875: sound1 <=  -386475;
	2876: sound1 <=  -312073;
	2877: sound1 <=  -245544;
	2878: sound1 <=  -148926;
	2879: sound1 <=  -56580;
	2880: sound1 <=  9064;
	2881: sound1 <=  90698;
	2882: sound1 <=  43945;
	2883: sound1 <=  -38635;
	2884: sound1 <=  -10925;
	2885: sound1 <=  8087;
	2886: sound1 <=  67688;
	2887: sound1 <=  100525;
	2888: sound1 <=  58655;
	2889: sound1 <=  -78918;
	2890: sound1 <=  -103119;
	2891: sound1 <=  -118958;
	2892: sound1 <=  -99243;
	2893: sound1 <=  -109100;
	2894: sound1 <=  -100098;
	2895: sound1 <=  -112579;
	2896: sound1 <=  -129913;
	2897: sound1 <=  -127899;
	2898: sound1 <=  -148010;
	2899: sound1 <=  -145599;
	2900: sound1 <=  -84137;
	2901: sound1 <=  -31586;
	2902: sound1 <=  24445;
	2903: sound1 <=  96008;
	2904: sound1 <=  143555;
	2905: sound1 <=  163879;
	2906: sound1 <=  187714;
	2907: sound1 <=  222717;
	2908: sound1 <=  277130;
	2909: sound1 <=  326599;
	2910: sound1 <=  353302;
	2911: sound1 <=  370880;
	2912: sound1 <=  378113;
	2913: sound1 <=  314392;
	2914: sound1 <=  279816;
	2915: sound1 <=  285767;
	2916: sound1 <=  313446;
	2917: sound1 <=  302429;
	2918: sound1 <=  316376;
	2919: sound1 <=  336121;
	2920: sound1 <=  326935;
	2921: sound1 <=  319092;
	2922: sound1 <=  322021;
	2923: sound1 <=  330566;
	2924: sound1 <=  333984;
	2925: sound1 <=  327148;
	2926: sound1 <=  316589;
	2927: sound1 <=  304504;
	2928: sound1 <=  316315;
	2929: sound1 <=  287048;
	2930: sound1 <=  266266;
	2931: sound1 <=  219330;
	2932: sound1 <=  137573;
	2933: sound1 <=  113098;
	2934: sound1 <=  128113;
	2935: sound1 <=  96252;
	2936: sound1 <=  56793;
	2937: sound1 <=  11139;
	2938: sound1 <=  -27069;
	2939: sound1 <=  -61005;
	2940: sound1 <=  -40314;
	2941: sound1 <=  -6104;
	2942: sound1 <=  -36316;
	2943: sound1 <=  -49835;
	2944: sound1 <=  -53955;
	2945: sound1 <=  -49500;
	2946: sound1 <=  -57831;
	2947: sound1 <=  -60211;
	2948: sound1 <=  -57434;
	2949: sound1 <=  -52551;
	2950: sound1 <=  -178772;
	2951: sound1 <=  -197784;
	2952: sound1 <=  -195465;
	2953: sound1 <=  -155090;
	2954: sound1 <=  -159668;
	2955: sound1 <=  -273254;
	2956: sound1 <=  -203339;
	2957: sound1 <=  -141846;
	2958: sound1 <=  -97107;
	2959: sound1 <=  -123596;
	2960: sound1 <=  -227142;
	2961: sound1 <=  -202026;
	2962: sound1 <=  -212250;
	2963: sound1 <=  -225677;
	2964: sound1 <=  -242920;
	2965: sound1 <=  -261566;
	2966: sound1 <=  -258514;
	2967: sound1 <=  -262207;
	2968: sound1 <=  -255707;
	2969: sound1 <=  -219177;
	2970: sound1 <=  -190155;
	2971: sound1 <=  -193390;
	2972: sound1 <=  -162231;
	2973: sound1 <=  -114685;
	2974: sound1 <=  -77454;
	2975: sound1 <=  -5829;
	2976: sound1 <=  51208;
	2977: sound1 <=  102753;
	2978: sound1 <=  107208;
	2979: sound1 <=  128326;
	2980: sound1 <=  101929;
	2981: sound1 <=  -33203;
	2982: sound1 <=  -50293;
	2983: sound1 <=  -85052;
	2984: sound1 <=  -40802;
	2985: sound1 <=  18005;
	2986: sound1 <=  43488;
	2987: sound1 <=  80383;
	2988: sound1 <=  122772;
	2989: sound1 <=  106079;
	2990: sound1 <=  -85754;
	2991: sound1 <=  -143951;
	2992: sound1 <=  -160065;
	2993: sound1 <=  -180878;
	2994: sound1 <=  -197571;
	2995: sound1 <=  -196381;
	2996: sound1 <=  -160736;
	2997: sound1 <=  -125122;
	2998: sound1 <=  -78430;
	2999: sound1 <=  -65247;
	3000: sound1 <=  -69061;
	3001: sound1 <=  -45959;
	3002: sound1 <=  5310;
	3003: sound1 <=  67810;
	3004: sound1 <=  116486;
	3005: sound1 <=  112885;
	3006: sound1 <=  169312;
	3007: sound1 <=  238800;
	3008: sound1 <=  256744;
	3009: sound1 <=  301208;
	3010: sound1 <=  326202;
	3011: sound1 <=  325958;
	3012: sound1 <=  330200;
	3013: sound1 <=  348206;
	3014: sound1 <=  365662;
	3015: sound1 <=  341309;
	3016: sound1 <=  338654;
	3017: sound1 <=  371704;
	3018: sound1 <=  404358;
	3019: sound1 <=  432648;
	3020: sound1 <=  416687;
	3021: sound1 <=  380829;
	3022: sound1 <=  344849;
	3023: sound1 <=  121155;
	3024: sound1 <=  -8301;
	3025: sound1 <=  -91644;
	3026: sound1 <=  -183777;
	3027: sound1 <=  -203461;
	3028: sound1 <=  -209412;
	3029: sound1 <=  -231232;
	3030: sound1 <=  -230896;
	3031: sound1 <=  -231598;
	3032: sound1 <=  -175201;
	3033: sound1 <=  -99915;
	3034: sound1 <=  -47119;
	3035: sound1 <=  13245;
	3036: sound1 <=  64026;
	3037: sound1 <=  121826;
	3038: sound1 <=  176514;
	3039: sound1 <=  160248;
	3040: sound1 <=  34607;
	3041: sound1 <=  41382;
	3042: sound1 <=  82275;
	3043: sound1 <=  136505;
	3044: sound1 <=  187592;
	3045: sound1 <=  138092;
	3046: sound1 <=  157135;
	3047: sound1 <=  181732;
	3048: sound1 <=  185394;
	3049: sound1 <=  116638;
	3050: sound1 <=  41473;
	3051: sound1 <=  125793;
	3052: sound1 <=  163788;
	3053: sound1 <=  79895;
	3054: sound1 <=  -54901;
	3055: sound1 <=  -83527;
	3056: sound1 <=  -82062;
	3057: sound1 <=  -41077;
	3058: sound1 <=  -30334;
	3059: sound1 <=  -31525;
	3060: sound1 <=  -34058;
	3061: sound1 <=  -119446;
	3062: sound1 <=  -145996;
	3063: sound1 <=  -131989;
	3064: sound1 <=  -155365;
	3065: sound1 <=  -159729;
	3066: sound1 <=  -146881;
	3067: sound1 <=  -126953;
	3068: sound1 <=  -121185;
	3069: sound1 <=  -116882;
	3070: sound1 <=  -93414;
	3071: sound1 <=  -84106;
	3072: sound1 <=  -57007;
	3073: sound1 <=  -20966;
	3074: sound1 <=  24719;
	3075: sound1 <=  60211;
	3076: sound1 <=  55817;
	3077: sound1 <=  95886;
	3078: sound1 <=  111298;
	3079: sound1 <=  96130;
	3080: sound1 <=  95215;
	3081: sound1 <=  86334;
	3082: sound1 <=  92133;
	3083: sound1 <=  86304;
	3084: sound1 <=  95978;
	3085: sound1 <=  111572;
	3086: sound1 <=  142853;
	3087: sound1 <=  198669;
	3088: sound1 <=  221069;
	3089: sound1 <=  220490;
	3090: sound1 <=  253082;
	3091: sound1 <=  309570;
	3092: sound1 <=  343628;
	3093: sound1 <=  319244;
	3094: sound1 <=  280243;
	3095: sound1 <=  263000;
	3096: sound1 <=  258423;
	3097: sound1 <=  270630;
	3098: sound1 <=  268921;
	3099: sound1 <=  253448;
	3100: sound1 <=  254120;
	3101: sound1 <=  296570;
	3102: sound1 <=  307678;
	3103: sound1 <=  303925;
	3104: sound1 <=  259827;
	3105: sound1 <=  199432;
	3106: sound1 <=  154907;
	3107: sound1 <=  92957;
	3108: sound1 <=  76874;
	3109: sound1 <=  57861;
	3110: sound1 <=  12543;
	3111: sound1 <=  -16998;
	3112: sound1 <=  -46082;
	3113: sound1 <=  -77881;
	3114: sound1 <=  -82825;
	3115: sound1 <=  -117615;
	3116: sound1 <=  -126160;
	3117: sound1 <=  -107849;
	3118: sound1 <=  -89752;
	3119: sound1 <=  -66376;
	3120: sound1 <=  -19989;
	3121: sound1 <=  18097;
	3122: sound1 <=  60547;
	3123: sound1 <=  69397;
	3124: sound1 <=  61981;
	3125: sound1 <=  81543;
	3126: sound1 <=  81390;
	3127: sound1 <=  72906;
	3128: sound1 <=  16998;
	3129: sound1 <=  -94421;
	3130: sound1 <=  -146790;
	3131: sound1 <=  -158600;
	3132: sound1 <=  -139618;
	3133: sound1 <=  -122742;
	3134: sound1 <=  -101410;
	3135: sound1 <=  -99426;
	3136: sound1 <=  -104218;
	3137: sound1 <=  -123840;
	3138: sound1 <=  -145081;
	3139: sound1 <=  -145294;
	3140: sound1 <=  -187378;
	3141: sound1 <=  -162781;
	3142: sound1 <=  -163544;
	3143: sound1 <=  -172089;
	3144: sound1 <=  -162201;
	3145: sound1 <=  -131165;
	3146: sound1 <=  -134369;
	3147: sound1 <=  -143066;
	3148: sound1 <=  -123047;
	3149: sound1 <=  -96161;
	3150: sound1 <=  -51666;
	3151: sound1 <=  -34363;
	3152: sound1 <=  -24658;
	3153: sound1 <=  -31494;
	3154: sound1 <=  -22705;
	3155: sound1 <=  -6317;
	3156: sound1 <=  17975;
	3157: sound1 <=  72937;
	3158: sound1 <=  120331;
	3159: sound1 <=  198547;
	3160: sound1 <=  246429;
	3161: sound1 <=  262726;
	3162: sound1 <=  285156;
	3163: sound1 <=  281494;
	3164: sound1 <=  288300;
	3165: sound1 <=  288605;
	3166: sound1 <=  298889;
	3167: sound1 <=  325012;
	3168: sound1 <=  336090;
	3169: sound1 <=  328156;
	3170: sound1 <=  302765;
	3171: sound1 <=  260895;
	3172: sound1 <=  196686;
	3173: sound1 <=  159851;
	3174: sound1 <=  141052;
	3175: sound1 <=  118927;
	3176: sound1 <=  98145;
	3177: sound1 <=  110626;
	3178: sound1 <=  -37384;
	3179: sound1 <=  -229858;
	3180: sound1 <=  -250885;
	3181: sound1 <=  -313965;
	3182: sound1 <=  -317688;
	3183: sound1 <=  -320129;
	3184: sound1 <=  -325714;
	3185: sound1 <=  -315491;
	3186: sound1 <=  -304749;
	3187: sound1 <=  -299744;
	3188: sound1 <=  -306061;
	3189: sound1 <=  -264557;
	3190: sound1 <=  -198151;
	3191: sound1 <=  -104004;
	3192: sound1 <=  -12970;
	3193: sound1 <=  66620;
	3194: sound1 <=  173004;
	3195: sound1 <=  236420;
	3196: sound1 <=  256897;
	3197: sound1 <=  327393;
	3198: sound1 <=  308044;
	3199: sound1 <=  300934;
	3200: sound1 <=  329773;
	3201: sound1 <=  342224;
	3202: sound1 <=  347198;
	3203: sound1 <=  299103;
	3204: sound1 <=  264252;
	3205: sound1 <=  318268;
	3206: sound1 <=  248077;
	3207: sound1 <=  196594;
	3208: sound1 <=  202728;
	3209: sound1 <=  206238;
	3210: sound1 <=  139343;
	3211: sound1 <=  60303;
	3212: sound1 <=  123810;
	3213: sound1 <=  29175;
	3214: sound1 <=  62744;
	3215: sound1 <=  -51239;
	3216: sound1 <=  -29663;
	3217: sound1 <=  -57373;
	3218: sound1 <=  -85724;
	3219: sound1 <=  -82031;
	3220: sound1 <=  -117798;
	3221: sound1 <=  -216431;
	3222: sound1 <=  -255463;
	3223: sound1 <=  -248474;
	3224: sound1 <=  -351746;
	3225: sound1 <=  -364838;
	3226: sound1 <=  -358307;
	3227: sound1 <=  -359497;
	3228: sound1 <=  -346436;
	3229: sound1 <=  -333038;
	3230: sound1 <=  -294006;
	3231: sound1 <=  -206726;
	3232: sound1 <=  -185791;
	3233: sound1 <=  -142181;
	3234: sound1 <=  -104126;
	3235: sound1 <=  -84412;
	3236: sound1 <=  -57190;
	3237: sound1 <=  -10864;
	3238: sound1 <=  -14984;
	3239: sound1 <=  -17334;
	3240: sound1 <=  -2991;
	3241: sound1 <=  1678;
	3242: sound1 <=  -18921;
	3243: sound1 <=  -33875;
	3244: sound1 <=  -99091;
	3245: sound1 <=  -46722;
	3246: sound1 <=  24719;
	3247: sound1 <=  -71259;
	3248: sound1 <=  -82458;
	3249: sound1 <=  -26489;
	3250: sound1 <=  40314;
	3251: sound1 <=  91461;
	3252: sound1 <=  148438;
	3253: sound1 <=  83496;
	3254: sound1 <=  -41443;
	3255: sound1 <=  25330;
	3256: sound1 <=  33081;
	3257: sound1 <=  39703;
	3258: sound1 <=  86548;
	3259: sound1 <=  21637;
	3260: sound1 <=  -96954;
	3261: sound1 <=  -71625;
	3262: sound1 <=  -3357;
	3263: sound1 <=  73059;
	3264: sound1 <=  143188;
	3265: sound1 <=  108337;
	3266: sound1 <=  47638;
	3267: sound1 <=  127106;
	3268: sound1 <=  152649;
	3269: sound1 <=  184204;
	3270: sound1 <=  95093;
	3271: sound1 <=  139374;
	3272: sound1 <=  192841;
	3273: sound1 <=  186096;
	3274: sound1 <=  120544;
	3275: sound1 <=  222778;
	3276: sound1 <=  319702;
	3277: sound1 <=  334167;
	3278: sound1 <=  258636;
	3279: sound1 <=  252686;
	3280: sound1 <=  216980;
	3281: sound1 <=  204041;
	3282: sound1 <=  215637;
	3283: sound1 <=  244354;
	3284: sound1 <=  291870;
	3285: sound1 <=  244171;
	3286: sound1 <=  158264;
	3287: sound1 <=  185181;
	3288: sound1 <=  130280;
	3289: sound1 <=  112183;
	3290: sound1 <=  108063;
	3291: sound1 <=  124115;
	3292: sound1 <=  156189;
	3293: sound1 <=  180176;
	3294: sound1 <=  44098;
	3295: sound1 <=  69611;
	3296: sound1 <=  128937;
	3297: sound1 <=  148468;
	3298: sound1 <=  73395;
	3299: sound1 <=  25116;
	3300: sound1 <=  79834;
	3301: sound1 <=  98785;
	3302: sound1 <=  97534;
	3303: sound1 <=  84106;
	3304: sound1 <=  56061;
	3305: sound1 <=  52643;
	3306: sound1 <=  51819;
	3307: sound1 <=  41840;
	3308: sound1 <=  83740;
	3309: sound1 <=  50354;
	3310: sound1 <=  -132446;
	3311: sound1 <=  -138153;
	3312: sound1 <=  -178711;
	3313: sound1 <=  -215240;
	3314: sound1 <=  -216888;
	3315: sound1 <=  -218414;
	3316: sound1 <=  -199738;
	3317: sound1 <=  -126984;
	3318: sound1 <=  -100861;
	3319: sound1 <=  -101105;
	3320: sound1 <=  -87585;
	3321: sound1 <=  -54535;
	3322: sound1 <=  -68939;
	3323: sound1 <=  -56854;
	3324: sound1 <=  21851;
	3325: sound1 <=  116638;
	3326: sound1 <=  215057;
	3327: sound1 <=  269714;
	3328: sound1 <=  298889;
	3329: sound1 <=  346436;
	3330: sound1 <=  380707;
	3331: sound1 <=  389648;
	3332: sound1 <=  390656;
	3333: sound1 <=  399933;
	3334: sound1 <=  377930;
	3335: sound1 <=  329712;
	3336: sound1 <=  299500;
	3337: sound1 <=  306152;
	3338: sound1 <=  299591;
	3339: sound1 <=  261719;
	3340: sound1 <=  229584;
	3341: sound1 <=  182495;
	3342: sound1 <=  144623;
	3343: sound1 <=  105438;
	3344: sound1 <=  53314;
	3345: sound1 <=  -75562;
	3346: sound1 <=  -308807;
	3347: sound1 <=  -383331;
	3348: sound1 <=  -450958;
	3349: sound1 <=  -498657;
	3350: sound1 <=  -501892;
	3351: sound1 <=  -506653;
	3352: sound1 <=  -496399;
	3353: sound1 <=  -474182;
	3354: sound1 <=  -450134;
	3355: sound1 <=  -451355;
	3356: sound1 <=  -442566;
	3357: sound1 <=  -426422;
	3358: sound1 <=  -399017;
	3359: sound1 <=  -389252;
	3360: sound1 <=  -371704;
	3361: sound1 <=  -303101;
	3362: sound1 <=  -221313;
	3363: sound1 <=  -154480;
	3364: sound1 <=  -94238;
	3365: sound1 <=  -59143;
	3366: sound1 <=  -36774;
	3367: sound1 <=  977;
	3368: sound1 <=  22400;
	3369: sound1 <=  33600;
	3370: sound1 <=  53284;
	3371: sound1 <=  59845;
	3372: sound1 <=  44250;
	3373: sound1 <=  73822;
	3374: sound1 <=  99213;
	3375: sound1 <=  96985;
	3376: sound1 <=  107239;
	3377: sound1 <=  113495;
	3378: sound1 <=  121033;
	3379: sound1 <=  107574;
	3380: sound1 <=  65582;
	3381: sound1 <=  22644;
	3382: sound1 <=  3387;
	3383: sound1 <=  -38544;
	3384: sound1 <=  -52002;
	3385: sound1 <=  -10956;
	3386: sound1 <=  13153;
	3387: sound1 <=  122;
	3388: sound1 <=  8087;
	3389: sound1 <=  -55328;
	3390: sound1 <=  -174408;
	3391: sound1 <=  -136292;
	3392: sound1 <=  -102325;
	3393: sound1 <=  -99091;
	3394: sound1 <=  -119446;
	3395: sound1 <=  -116425;
	3396: sound1 <=  -109894;
	3397: sound1 <=  -90515;
	3398: sound1 <=  -77301;
	3399: sound1 <=  -81177;
	3400: sound1 <=  -77148;
	3401: sound1 <=  -60547;
	3402: sound1 <=  -38177;
	3403: sound1 <=  -22675;
	3404: sound1 <=  11597;
	3405: sound1 <=  56763;
	3406: sound1 <=  117889;
	3407: sound1 <=  169556;
	3408: sound1 <=  287262;
	3409: sound1 <=  387787;
	3410: sound1 <=  414154;
	3411: sound1 <=  451935;
	3412: sound1 <=  478882;
	3413: sound1 <=  506500;
	3414: sound1 <=  549988;
	3415: sound1 <=  582581;
	3416: sound1 <=  614899;
	3417: sound1 <=  635681;
	3418: sound1 <=  633820;
	3419: sound1 <=  581573;
	3420: sound1 <=  529968;
	3421: sound1 <=  507751;
	3422: sound1 <=  455963;
	3423: sound1 <=  425385;
	3424: sound1 <=  406647;
	3425: sound1 <=  381592;
	3426: sound1 <=  359772;
	3427: sound1 <=  328644;
	3428: sound1 <=  276703;
	3429: sound1 <=  238678;
	3430: sound1 <=  194153;
	3431: sound1 <=  113373;
	3432: sound1 <=  40131;
	3433: sound1 <=  28717;
	3434: sound1 <=  -5798;
	3435: sound1 <=  -60699;
	3436: sound1 <=  -132660;
	3437: sound1 <=  -181763;
	3438: sound1 <=  -198395;
	3439: sound1 <=  -207947;
	3440: sound1 <=  -215546;
	3441: sound1 <=  -186584;
	3442: sound1 <=  -160187;
	3443: sound1 <=  -156616;
	3444: sound1 <=  -151611;
	3445: sound1 <=  -157745;
	3446: sound1 <=  -153839;
	3447: sound1 <=  -160522;
	3448: sound1 <=  -175110;
	3449: sound1 <=  -160797;
	3450: sound1 <=  -122711;
	3451: sound1 <=  -108521;
	3452: sound1 <=  -127258;
	3453: sound1 <=  -152771;
	3454: sound1 <=  -172729;
	3455: sound1 <=  -145233;
	3456: sound1 <=  -128876;
	3457: sound1 <=  -66711;
	3458: sound1 <=  -42450;
	3459: sound1 <=  -54169;
	3460: sound1 <=  -72235;
	3461: sound1 <=  -100403;
	3462: sound1 <=  -132355;
	3463: sound1 <=  -169769;
	3464: sound1 <=  -207947;
	3465: sound1 <=  -241730;
	3466: sound1 <=  -218231;
	3467: sound1 <=  -195709;
	3468: sound1 <=  -220001;
	3469: sound1 <=  -236664;
	3470: sound1 <=  -231659;
	3471: sound1 <=  -235901;
	3472: sound1 <=  -225128;
	3473: sound1 <=  -208588;
	3474: sound1 <=  -191101;
	3475: sound1 <=  -184265;
	3476: sound1 <=  -216919;
	3477: sound1 <=  -243347;
	3478: sound1 <=  -266357;
	3479: sound1 <=  -279663;
	3480: sound1 <=  -266602;
	3481: sound1 <=  -255554;
	3482: sound1 <=  -263184;
	3483: sound1 <=  -258087;
	3484: sound1 <=  -227142;
	3485: sound1 <=  -201996;
	3486: sound1 <=  -158813;
	3487: sound1 <=  -157288;
	3488: sound1 <=  -165588;
	3489: sound1 <=  -165405;
	3490: sound1 <=  -166901;
	3491: sound1 <=  -136230;
	3492: sound1 <=  -101746;
	3493: sound1 <=  -102905;
	3494: sound1 <=  -104950;
	3495: sound1 <=  -88348;
	3496: sound1 <=  -16449;
	3497: sound1 <=  50323;
	3498: sound1 <=  89844;
	3499: sound1 <=  172028;
	3500: sound1 <=  278259;
	3501: sound1 <=  388397;
	3502: sound1 <=  482819;
	3503: sound1 <=  561615;
	3504: sound1 <=  649780;
	3505: sound1 <=  690460;
	3506: sound1 <=  727692;
	3507: sound1 <=  747925;
	3508: sound1 <=  764435;
	3509: sound1 <=  742340;
	3510: sound1 <=  695190;
	3511: sound1 <=  625488;
	3512: sound1 <=  575623;
	3513: sound1 <=  545013;
	3514: sound1 <=  523102;
	3515: sound1 <=  443512;
	3516: sound1 <=  351044;
	3517: sound1 <=  305664;
	3518: sound1 <=  296417;
	3519: sound1 <=  265320;
	3520: sound1 <=  220184;
	3521: sound1 <=  173889;
	3522: sound1 <=  129425;
	3523: sound1 <=  98694;
	3524: sound1 <=  106873;
	3525: sound1 <=  127441;
	3526: sound1 <=  132202;
	3527: sound1 <=  121429;
	3528: sound1 <=  107086;
	3529: sound1 <=  98175;
	3530: sound1 <=  101929;
	3531: sound1 <=  113892;
	3532: sound1 <=  83008;
	3533: sound1 <=  53162;
	3534: sound1 <=  37201;
	3535: sound1 <=  -19989;
	3536: sound1 <=  -60974;
	3537: sound1 <=  -73975;
	3538: sound1 <=  -73273;
	3539: sound1 <=  -82642;
	3540: sound1 <=  -97198;
	3541: sound1 <=  -97382;
	3542: sound1 <=  -238190;
	3543: sound1 <=  -329498;
	3544: sound1 <=  -299133;
	3545: sound1 <=  -303558;
	3546: sound1 <=  -295898;
	3547: sound1 <=  -317596;
	3548: sound1 <=  -317139;
	3549: sound1 <=  -315552;
	3550: sound1 <=  -285889;
	3551: sound1 <=  -295288;
	3552: sound1 <=  -285553;
	3553: sound1 <=  -256409;
	3554: sound1 <=  -219940;
	3555: sound1 <=  -156494;
	3556: sound1 <=  -69061;
	3557: sound1 <=  25696;
	3558: sound1 <=  83038;
	3559: sound1 <=  105255;
	3560: sound1 <=  133881;
	3561: sound1 <=  196747;
	3562: sound1 <=  219574;
	3563: sound1 <=  208099;
	3564: sound1 <=  192749;
	3565: sound1 <=  11963;
	3566: sound1 <=  -133484;
	3567: sound1 <=  -121887;
	3568: sound1 <=  -125610;
	3569: sound1 <=  -127594;
	3570: sound1 <=  -133606;
	3571: sound1 <=  -115234;
	3572: sound1 <=  -103119;
	3573: sound1 <=  -96710;
	3574: sound1 <=  -84808;
	3575: sound1 <=  -89569;
	3576: sound1 <=  -109924;
	3577: sound1 <=  -147003;
	3578: sound1 <=  -150574;
	3579: sound1 <=  -116638;
	3580: sound1 <=  -86304;
	3581: sound1 <=  -14526;
	3582: sound1 <=  73639;
	3583: sound1 <=  125153;
	3584: sound1 <=  188202;
	3585: sound1 <=  241608;
	3586: sound1 <=  293976;
	3587: sound1 <=  324280;
	3588: sound1 <=  344910;
	3589: sound1 <=  373901;
	3590: sound1 <=  402649;
	3591: sound1 <=  405457;
	3592: sound1 <=  400269;
	3593: sound1 <=  415253;
	3594: sound1 <=  436432;
	3595: sound1 <=  446899;
	3596: sound1 <=  449371;
	3597: sound1 <=  437378;
	3598: sound1 <=  383728;
	3599: sound1 <=  336578;
	3600: sound1 <=  308319;
	3601: sound1 <=  264893;
	3602: sound1 <=  231018;
	3603: sound1 <=  201874;
	3604: sound1 <=  162262;
	3605: sound1 <=  79315;
	3606: sound1 <=  39673;
	3607: sound1 <=  -147308;
	3608: sound1 <=  -267303;
	3609: sound1 <=  -304199;
	3610: sound1 <=  -345581;
	3611: sound1 <=  -358002;
	3612: sound1 <=  -398987;
	3613: sound1 <=  -429382;
	3614: sound1 <=  -430267;
	3615: sound1 <=  -423065;
	3616: sound1 <=  -393005;
	3617: sound1 <=  -309692;
	3618: sound1 <=  -253479;
	3619: sound1 <=  -254303;
	3620: sound1 <=  -229675;
	3621: sound1 <=  -214630;
	3622: sound1 <=  -173645;
	3623: sound1 <=  -107941;
	3624: sound1 <=  -66956;
	3625: sound1 <=  -4272;
	3626: sound1 <=  85083;
	3627: sound1 <=  70892;
	3628: sound1 <=  -30396;
	3629: sound1 <=  -28015;
	3630: sound1 <=  -46936;
	3631: sound1 <=  -32043;
	3632: sound1 <=  23865;
	3633: sound1 <=  67535;
	3634: sound1 <=  88257;
	3635: sound1 <=  85663;
	3636: sound1 <=  103455;
	3637: sound1 <=  103577;
	3638: sound1 <=  102539;
	3639: sound1 <=  -36011;
	3640: sound1 <=  -95703;
	3641: sound1 <=  -112488;
	3642: sound1 <=  -141815;
	3643: sound1 <=  -147247;
	3644: sound1 <=  -134949;
	3645: sound1 <=  -122131;
	3646: sound1 <=  -113617;
	3647: sound1 <=  -130157;
	3648: sound1 <=  -163055;
	3649: sound1 <=  -146088;
	3650: sound1 <=  -98328;
	3651: sound1 <=  -78583;
	3652: sound1 <=  -63324;
	3653: sound1 <=  -54932;
	3654: sound1 <=  -32684;
	3655: sound1 <=  14679;
	3656: sound1 <=  40771;
	3657: sound1 <=  105560;
	3658: sound1 <=  175812;
	3659: sound1 <=  202484;
	3660: sound1 <=  181946;
	3661: sound1 <=  175812;
	3662: sound1 <=  213196;
	3663: sound1 <=  216156;
	3664: sound1 <=  223145;
	3665: sound1 <=  274902;
	3666: sound1 <=  331573;
	3667: sound1 <=  383514;
	3668: sound1 <=  423035;
	3669: sound1 <=  443542;
	3670: sound1 <=  460419;
	3671: sound1 <=  454559;
	3672: sound1 <=  462921;
	3673: sound1 <=  439301;
	3674: sound1 <=  388824;
	3675: sound1 <=  339111;
	3676: sound1 <=  283600;
	3677: sound1 <=  238586;
	3678: sound1 <=  190887;
	3679: sound1 <=  222870;
	3680: sound1 <=  248108;
	3681: sound1 <=  228424;
	3682: sound1 <=  219757;
	3683: sound1 <=  218140;
	3684: sound1 <=  187195;
	3685: sound1 <=  133545;
	3686: sound1 <=  83099;
	3687: sound1 <=  28320;
	3688: sound1 <=  -8423;
	3689: sound1 <=  -66345;
	3690: sound1 <=  -69000;
	3691: sound1 <=  -48004;
	3692: sound1 <=  -44678;
	3693: sound1 <=  -74036;
	3694: sound1 <=  -103546;
	3695: sound1 <=  -97504;
	3696: sound1 <=  -87067;
	3697: sound1 <=  -63995;
	3698: sound1 <=  -45410;
	3699: sound1 <=  -61493;
	3700: sound1 <=  -47699;
	3701: sound1 <=  -3571;
	3702: sound1 <=  1648;
	3703: sound1 <=  -3723;
	3704: sound1 <=  -2197;
	3705: sound1 <=  13550;
	3706: sound1 <=  5341;
	3707: sound1 <=  -13550;
	3708: sound1 <=  -41046;
	3709: sound1 <=  -90698;
	3710: sound1 <=  -157776;
	3711: sound1 <=  -184875;
	3712: sound1 <=  -200165;
	3713: sound1 <=  -230347;
	3714: sound1 <=  -250214;
	3715: sound1 <=  -256104;
	3716: sound1 <=  -216827;
	3717: sound1 <=  -226227;
	3718: sound1 <=  -269135;
	3719: sound1 <=  -333801;
	3720: sound1 <=  -341461;
	3721: sound1 <=  -321503;
	3722: sound1 <=  -331848;
	3723: sound1 <=  -288086;
	3724: sound1 <=  -255371;
	3725: sound1 <=  -197693;
	3726: sound1 <=  -142487;
	3727: sound1 <=  -78125;
	3728: sound1 <=  -75378;
	3729: sound1 <=  -68329;
	3730: sound1 <=  -58014;
	3731: sound1 <=  -58502;
	3732: sound1 <=  -13824;
	3733: sound1 <=  16632;
	3734: sound1 <=  -18829;
	3735: sound1 <=  -56427;
	3736: sound1 <=  -74829;
	3737: sound1 <=  -57159;
	3738: sound1 <=  -63965;
	3739: sound1 <=  -59204;
	3740: sound1 <=  -41748;
	3741: sound1 <=  -18921;
	3742: sound1 <=  -7080;
	3743: sound1 <=  -44525;
	3744: sound1 <=  -50568;
	3745: sound1 <=  -55573;
	3746: sound1 <=  -147217;
	3747: sound1 <=  -120300;
	3748: sound1 <=  -92316;
	3749: sound1 <=  -75348;
	3750: sound1 <=  -73761;
	3751: sound1 <=  -76813;
	3752: sound1 <=  -101837;
	3753: sound1 <=  -118317;
	3754: sound1 <=  -120636;
	3755: sound1 <=  -104736;
	3756: sound1 <=  -69458;
	3757: sound1 <=  -47699;
	3758: sound1 <=  -14679;
	3759: sound1 <=  30579;
	3760: sound1 <=  53589;
	3761: sound1 <=  87402;
	3762: sound1 <=  159271;
	3763: sound1 <=  219055;
	3764: sound1 <=  243774;
	3765: sound1 <=  306488;
	3766: sound1 <=  313110;
	3767: sound1 <=  321655;
	3768: sound1 <=  316193;
	3769: sound1 <=  302521;
	3770: sound1 <=  312134;
	3771: sound1 <=  339630;
	3772: sound1 <=  334747;
	3773: sound1 <=  348053;
	3774: sound1 <=  359314;
	3775: sound1 <=  387054;
	3776: sound1 <=  402313;
	3777: sound1 <=  402313;
	3778: sound1 <=  408386;
	3779: sound1 <=  400879;
	3780: sound1 <=  384308;
	3781: sound1 <=  354004;
	3782: sound1 <=  347260;
	3783: sound1 <=  239990;
	3784: sound1 <=  129028;
	3785: sound1 <=  161804;
	3786: sound1 <=  158936;
	3787: sound1 <=  140167;
	3788: sound1 <=  123657;
	3789: sound1 <=  128143;
	3790: sound1 <=  114990;
	3791: sound1 <=  81909;
	3792: sound1 <=  28992;
	3793: sound1 <=  8301;
	3794: sound1 <=  2441;
	3795: sound1 <=  519;
	3796: sound1 <=  -4303;
	3797: sound1 <=  21667;
	3798: sound1 <=  51636;
	3799: sound1 <=  32501;
	3800: sound1 <=  33112;
	3801: sound1 <=  32410;
	3802: sound1 <=  92;
	3803: sound1 <=  -20844;
	3804: sound1 <=  -32501;
	3805: sound1 <=  -189453;
	3806: sound1 <=  -299957;
	3807: sound1 <=  -377655;
	3808: sound1 <=  -384094;
	3809: sound1 <=  -373230;
	3810: sound1 <=  -372681;
	3811: sound1 <=  -330170;
	3812: sound1 <=  -280457;
	3813: sound1 <=  -238007;
	3814: sound1 <=  -166870;
	3815: sound1 <=  -72601;
	3816: sound1 <=  18280;
	3817: sound1 <=  98511;
	3818: sound1 <=  76324;
	3819: sound1 <=  12634;
	3820: sound1 <=  83130;
	3821: sound1 <=  124146;
	3822: sound1 <=  185852;
	3823: sound1 <=  222717;
	3824: sound1 <=  229431;
	3825: sound1 <=  95245;
	3826: sound1 <=  60364;
	3827: sound1 <=  63965;
	3828: sound1 <=  44983;
	3829: sound1 <=  33875;
	3830: sound1 <=  16907;
	3831: sound1 <=  3204;
	3832: sound1 <=  -3906;
	3833: sound1 <=  12421;
	3834: sound1 <=  43884;
	3835: sound1 <=  69458;
	3836: sound1 <=  66345;
	3837: sound1 <=  73975;
	3838: sound1 <=  82428;
	3839: sound1 <=  62683;
	3840: sound1 <=  -11383;
	3841: sound1 <=  -152679;
	3842: sound1 <=  -160126;
	3843: sound1 <=  -167908;
	3844: sound1 <=  -173615;
	3845: sound1 <=  -153259;
	3846: sound1 <=  -141052;
	3847: sound1 <=  -142181;
	3848: sound1 <=  -160736;
	3849: sound1 <=  -164215;
	3850: sound1 <=  -152802;
	3851: sound1 <=  -123444;
	3852: sound1 <=  -89813;
	3853: sound1 <=  -33356;
	3854: sound1 <=  35767;
	3855: sound1 <=  65674;
	3856: sound1 <=  113586;
	3857: sound1 <=  193329;
	3858: sound1 <=  250824;
	3859: sound1 <=  274536;
	3860: sound1 <=  265198;
	3861: sound1 <=  305450;
	3862: sound1 <=  360382;
	3863: sound1 <=  394073;
	3864: sound1 <=  399902;
	3865: sound1 <=  420044;
	3866: sound1 <=  418549;
	3867: sound1 <=  402557;
	3868: sound1 <=  367737;
	3869: sound1 <=  339264;
	3870: sound1 <=  332642;
	3871: sound1 <=  339996;
	3872: sound1 <=  308197;
	3873: sound1 <=  286865;
	3874: sound1 <=  263123;
	3875: sound1 <=  186737;
	3876: sound1 <=  145172;
	3877: sound1 <=  79437;
	3878: sound1 <=  -135590;
	3879: sound1 <=  -157410;
	3880: sound1 <=  -184601;
	3881: sound1 <=  -207184;
	3882: sound1 <=  -200348;
	3883: sound1 <=  -191986;
	3884: sound1 <=  -160370;
	3885: sound1 <=  -122131;
	3886: sound1 <=  -90332;
	3887: sound1 <=  -68268;
	3888: sound1 <=  -67078;
	3889: sound1 <=  -46936;
	3890: sound1 <=  -5463;
	3891: sound1 <=  31464;
	3892: sound1 <=  70892;
	3893: sound1 <=  -52307;
	3894: sound1 <=  -122620;
	3895: sound1 <=  -112579;
	3896: sound1 <=  -125000;
	3897: sound1 <=  -158142;
	3898: sound1 <=  -176117;
	3899: sound1 <=  -158936;
	3900: sound1 <=  -155731;
	3901: sound1 <=  -142822;
	3902: sound1 <=  -113525;
	3903: sound1 <=  -92072;
	3904: sound1 <=  -109161;
	3905: sound1 <=  -72845;
	3906: sound1 <=  -71747;
	3907: sound1 <=  -72968;
	3908: sound1 <=  -149414;
	3909: sound1 <=  -283203;
	3910: sound1 <=  -242401;
	3911: sound1 <=  -232361;
	3912: sound1 <=  -222321;
	3913: sound1 <=  -204803;
	3914: sound1 <=  -199677;
	3915: sound1 <=  -179932;
	3916: sound1 <=  -149414;
	3917: sound1 <=  -130920;
	3918: sound1 <=  -128876;
	3919: sound1 <=  -94757;
	3920: sound1 <=  -12787;
	3921: sound1 <=  102051;
	3922: sound1 <=  187164;
	3923: sound1 <=  259338;
	3924: sound1 <=  318665;
	3925: sound1 <=  340790;
	3926: sound1 <=  367737;
	3927: sound1 <=  358704;
	3928: sound1 <=  329010;
	3929: sound1 <=  344940;
	3930: sound1 <=  353180;
	3931: sound1 <=  354950;
	3932: sound1 <=  403748;
	3933: sound1 <=  452545;
	3934: sound1 <=  456421;
	3935: sound1 <=  436462;
	3936: sound1 <=  411255;
	3937: sound1 <=  423309;
	3938: sound1 <=  312042;
	3939: sound1 <=  113434;
	3940: sound1 <=  13245;
	3941: sound1 <=  -81818;
	3942: sound1 <=  -119781;
	3943: sound1 <=  -191315;
	3944: sound1 <=  -227570;
	3945: sound1 <=  -246796;
	3946: sound1 <=  -303528;
	3947: sound1 <=  -327759;
	3948: sound1 <=  -324188;
	3949: sound1 <=  -304047;
	3950: sound1 <=  -279327;
	3951: sound1 <=  -278809;
	3952: sound1 <=  -254486;
	3953: sound1 <=  -191071;
	3954: sound1 <=  -144989;
	3955: sound1 <=  -124268;
	3956: sound1 <=  -80200;
	3957: sound1 <=  -23956;
	3958: sound1 <=  13641;
	3959: sound1 <=  49683;
	3960: sound1 <=  99487;
	3961: sound1 <=  149902;
	3962: sound1 <=  158112;
	3963: sound1 <=  191223;
	3964: sound1 <=  186066;
	3965: sound1 <=  212952;
	3966: sound1 <=  247528;
	3967: sound1 <=  268768;
	3968: sound1 <=  277374;
	3969: sound1 <=  274261;
	3970: sound1 <=  258087;
	3971: sound1 <=  235016;
	3972: sound1 <=  195282;
	3973: sound1 <=  167053;
	3974: sound1 <=  161713;
	3975: sound1 <=  135712;
	3976: sound1 <=  136017;
	3977: sound1 <=  120209;
	3978: sound1 <=  103241;
	3979: sound1 <=  102448;
	3980: sound1 <=  75897;
	3981: sound1 <=  69824;
	3982: sound1 <=  29236;
	3983: sound1 <=  30121;
	3984: sound1 <=  10284;
	3985: sound1 <=  16907;
	3986: sound1 <=  18890;
	3987: sound1 <=  -5463;
	3988: sound1 <=  -32867;
	3989: sound1 <=  -36621;
	3990: sound1 <=  -23254;
	3991: sound1 <=  -12634;
	3992: sound1 <=  -28595;
	3993: sound1 <=  -38879;
	3994: sound1 <=  -50690;
	3995: sound1 <=  -46875;
	3996: sound1 <=  -44556;
	3997: sound1 <=  -72449;
	3998: sound1 <=  -129333;
	3999: sound1 <=  -138855;
	4000: sound1 <=  -104828;
	4001: sound1 <=  -95032;
	4002: sound1 <=  -106201;
	4003: sound1 <=  -105347;
	4004: sound1 <=  -106598;
	4005: sound1 <=  -83954;
	4006: sound1 <=  -65460;
	4007: sound1 <=  -43549;
	4008: sound1 <=  -45410;
	4009: sound1 <=  -37292;
	4010: sound1 <=  -5737;
	4011: sound1 <=  -18677;
	4012: sound1 <=  -50934;
	4013: sound1 <=  -58167;
	4014: sound1 <=  -64697;
	4015: sound1 <=  -50385;
	4016: sound1 <=  -43396;
	4017: sound1 <=  -46173;
	4018: sound1 <=  -75043;
	4019: sound1 <=  -97656;
	4020: sound1 <=  -89569;
	4021: sound1 <=  -81726;
	4022: sound1 <=  -40466;
	4023: sound1 <=  -16205;
	4024: sound1 <=  -11261;
	4025: sound1 <=  -14862;
	4026: sound1 <=  -1923;
	4027: sound1 <=  23529;
	4028: sound1 <=  27405;
	4029: sound1 <=  25726;
	4030: sound1 <=  13275;
	4031: sound1 <=  5310;
	4032: sound1 <=  -18829;
	4033: sound1 <=  -31769;
	4034: sound1 <=  -43762;
	4035: sound1 <=  -14984;
	4036: sound1 <=  16632;
	4037: sound1 <=  33447;
	4038: sound1 <=  70038;
	4039: sound1 <=  88623;
	4040: sound1 <=  99640;
	4041: sound1 <=  91125;
	4042: sound1 <=  70313;
	4043: sound1 <=  67902;
	4044: sound1 <=  68146;
	4045: sound1 <=  38055;
	4046: sound1 <=  47577;
	4047: sound1 <=  66986;
	4048: sound1 <=  96252;
	4049: sound1 <=  96954;
	4050: sound1 <=  70679;
	4051: sound1 <=  67169;
	4052: sound1 <=  83801;
	4053: sound1 <=  92072;
	4054: sound1 <=  102295;
	4055: sound1 <=  96741;
	4056: sound1 <=  -61646;
	4057: sound1 <=  -114838;
	4058: sound1 <=  -122192;
	4059: sound1 <=  -159546;
	4060: sound1 <=  -170776;
	4061: sound1 <=  -165131;
	4062: sound1 <=  -170685;
	4063: sound1 <=  -197479;
	4064: sound1 <=  -179962;
	4065: sound1 <=  -149200;
	4066: sound1 <=  -116852;
	4067: sound1 <=  -85266;
	4068: sound1 <=  -68268;
	4069: sound1 <=  -38300;
	4070: sound1 <=  1617;
	4071: sound1 <=  13275;
	4072: sound1 <=  24384;
	4073: sound1 <=  47150;
	4074: sound1 <=  77332;
	4075: sound1 <=  142456;
	4076: sound1 <=  214447;
	4077: sound1 <=  279785;
	4078: sound1 <=  323792;
	4079: sound1 <=  331665;
	4080: sound1 <=  340240;
	4081: sound1 <=  351227;
	4082: sound1 <=  333435;
	4083: sound1 <=  321838;
	4084: sound1 <=  347748;
	4085: sound1 <=  369019;
	4086: sound1 <=  388367;
	4087: sound1 <=  402100;
	4088: sound1 <=  411591;
	4089: sound1 <=  415009;
	4090: sound1 <=  429688;
	4091: sound1 <=  434723;
	4092: sound1 <=  432648;
	4093: sound1 <=  406952;
	4094: sound1 <=  346283;
	4095: sound1 <=  306305;
	4096: sound1 <=  292297;
	4097: sound1 <=  256073;
	4098: sound1 <=  214783;
	4099: sound1 <=  206787;
	4100: sound1 <=  200562;
	4101: sound1 <=  212158;
	4102: sound1 <=  205719;
	4103: sound1 <=  193420;
	4104: sound1 <=  193939;
	4105: sound1 <=  190399;
	4106: sound1 <=  177979;
	4107: sound1 <=  153046;
	4108: sound1 <=  146088;
	4109: sound1 <=  118988;
	4110: sound1 <=  98236;
	4111: sound1 <=  64026;
	4112: sound1 <=  42084;
	4113: sound1 <=  40039;
	4114: sound1 <=  15686;
	4115: sound1 <=  -19684;
	4116: sound1 <=  -78491;
	4117: sound1 <=  -111908;
	4118: sound1 <=  -121582;
	4119: sound1 <=  -139435;
	4120: sound1 <=  -155212;
	4121: sound1 <=  -150665;
	4122: sound1 <=  -162506;
	4123: sound1 <=  -157837;
	4124: sound1 <=  -153259;
	4125: sound1 <=  -178955;
	4126: sound1 <=  -265869;
	4127: sound1 <=  -282867;
	4128: sound1 <=  -266052;
	4129: sound1 <=  -298615;
	4130: sound1 <=  -339935;
	4131: sound1 <=  -372620;
	4132: sound1 <=  -401550;
	4133: sound1 <=  -388428;
	4134: sound1 <=  -378601;
	4135: sound1 <=  -391907;
	4136: sound1 <=  -392792;
	4137: sound1 <=  -370087;
	4138: sound1 <=  -329468;
	4139: sound1 <=  -301361;
	4140: sound1 <=  -273468;
	4141: sound1 <=  -228943;
	4142: sound1 <=  -213379;
	4143: sound1 <=  -171967;
	4144: sound1 <=  -83160;
	4145: sound1 <=  5432;
	4146: sound1 <=  73486;
	4147: sound1 <=  130310;
	4148: sound1 <=  151276;
	4149: sound1 <=  173859;
	4150: sound1 <=  194946;
	4151: sound1 <=  228668;
	4152: sound1 <=  283264;
	4153: sound1 <=  320129;
	4154: sound1 <=  336792;
	4155: sound1 <=  350098;
	4156: sound1 <=  328613;
	4157: sound1 <=  268829;
	4158: sound1 <=  232971;
	4159: sound1 <=  223389;
	4160: sound1 <=  206268;
	4161: sound1 <=  193787;
	4162: sound1 <=  187408;
	4163: sound1 <=  155701;
	4164: sound1 <=  146790;
	4165: sound1 <=  133545;
	4166: sound1 <=  107422;
	4167: sound1 <=  103241;
	4168: sound1 <=  94238;
	4169: sound1 <=  40894;
	4170: sound1 <=  12573;
	4171: sound1 <=  24841;
	4172: sound1 <=  9918;
	4173: sound1 <=  5280;
	4174: sound1 <=  22064;
	4175: sound1 <=  25940;
	4176: sound1 <=  2441;
	4177: sound1 <=  -21759;
	4178: sound1 <=  946;
	4179: sound1 <=  7996;
	4180: sound1 <=  -6561;
	4181: sound1 <=  -36652;
	4182: sound1 <=  -73730;
	4183: sound1 <=  -58624;
	4184: sound1 <=  -13489;
	4185: sound1 <=  -1617;
	4186: sound1 <=  -5981;
	4187: sound1 <=  6287;
	4188: sound1 <=  38727;
	4189: sound1 <=  48401;
	4190: sound1 <=  65460;
	4191: sound1 <=  81665;
	4192: sound1 <=  55206;
	4193: sound1 <=  28717;
	4194: sound1 <=  16479;
	4195: sound1 <=  -4761;
	4196: sound1 <=  -48279;
	4197: sound1 <=  -209076;
	4198: sound1 <=  -225800;
	4199: sound1 <=  -228241;
	4200: sound1 <=  -216309;
	4201: sound1 <=  -202728;
	4202: sound1 <=  -221832;
	4203: sound1 <=  -243622;
	4204: sound1 <=  -258026;
	4205: sound1 <=  -289795;
	4206: sound1 <=  -322418;
	4207: sound1 <=  -336517;
	4208: sound1 <=  -344299;
	4209: sound1 <=  -285431;
	4210: sound1 <=  -251526;
	4211: sound1 <=  -195465;
	4212: sound1 <=  -109863;
	4213: sound1 <=  -72784;
	4214: sound1 <=  -6409;
	4215: sound1 <=  47577;
	4216: sound1 <=  66956;
	4217: sound1 <=  87646;
	4218: sound1 <=  113281;
	4219: sound1 <=  177490;
	4220: sound1 <=  240753;
	4221: sound1 <=  284485;
	4222: sound1 <=  331360;
	4223: sound1 <=  378998;
	4224: sound1 <=  415955;
	4225: sound1 <=  421143;
	4226: sound1 <=  432312;
	4227: sound1 <=  413300;
	4228: sound1 <=  373749;
	4229: sound1 <=  330994;
	4230: sound1 <=  337036;
	4231: sound1 <=  349243;
	4232: sound1 <=  350006;
	4233: sound1 <=  345825;
	4234: sound1 <=  330933;
	4235: sound1 <=  308411;
	4236: sound1 <=  256012;
	4237: sound1 <=  192810;
	4238: sound1 <=  131134;
	4239: sound1 <=  99274;
	4240: sound1 <=  54901;
	4241: sound1 <=  23346;
	4242: sound1 <=  22186;
	4243: sound1 <=  35339;
	4244: sound1 <=  34393;
	4245: sound1 <=  20844;
	4246: sound1 <=  17242;
	4247: sound1 <=  8850;
	4248: sound1 <=  15900;
	4249: sound1 <=  22186;
	4250: sound1 <=  26947;
	4251: sound1 <=  25787;
	4252: sound1 <=  -3937;
	4253: sound1 <=  -31372;
	4254: sound1 <=  -82123;
	4255: sound1 <=  -123962;
	4256: sound1 <=  -147644;
	4257: sound1 <=  -160797;
	4258: sound1 <=  -171234;
	4259: sound1 <=  -206909;
	4260: sound1 <=  -239899;
	4261: sound1 <=  -261871;
	4262: sound1 <=  -248199;
	4263: sound1 <=  -244843;
	4264: sound1 <=  -264679;
	4265: sound1 <=  -290131;
	4266: sound1 <=  -289032;
	4267: sound1 <=  -267151;
	4268: sound1 <=  -237366;
	4269: sound1 <=  -220337;
	4270: sound1 <=  -243195;
	4271: sound1 <=  -260406;
	4272: sound1 <=  -246338;
	4273: sound1 <=  -214935;
	4274: sound1 <=  -187653;
	4275: sound1 <=  -175201;
	4276: sound1 <=  -179565;
	4277: sound1 <=  -178894;
	4278: sound1 <=  -162415;
	4279: sound1 <=  -123749;
	4280: sound1 <=  -66833;
	4281: sound1 <=  -75012;
	4282: sound1 <=  -70679;
	4283: sound1 <=  -67719;
	4284: sound1 <=  -75684;
	4285: sound1 <=  -78247;
	4286: sound1 <=  -68237;
	4287: sound1 <=  -37659;
	4288: sound1 <=  -18005;
	4289: sound1 <=  -885;
	4290: sound1 <=  3815;
	4291: sound1 <=  -15076;
	4292: sound1 <=  5371;
	4293: sound1 <=  91309;
	4294: sound1 <=  139191;
	4295: sound1 <=  184540;
	4296: sound1 <=  210815;
	4297: sound1 <=  213409;
	4298: sound1 <=  196716;
	4299: sound1 <=  204987;
	4300: sound1 <=  198578;
	4301: sound1 <=  199707;
	4302: sound1 <=  207062;
	4303: sound1 <=  204285;
	4304: sound1 <=  224030;
	4305: sound1 <=  266998;
	4306: sound1 <=  301331;
	4307: sound1 <=  278442;
	4308: sound1 <=  255646;
	4309: sound1 <=  144806;
	4310: sound1 <=  26642;
	4311: sound1 <=  18677;
	4312: sound1 <=  -32349;
	4313: sound1 <=  -42053;
	4314: sound1 <=  -82397;
	4315: sound1 <=  -94116;
	4316: sound1 <=  -82672;
	4317: sound1 <=  -82642;
	4318: sound1 <=  -88257;
	4319: sound1 <=  -51270;
	4320: sound1 <=  -20325;
	4321: sound1 <=  24292;
	4322: sound1 <=  65948;
	4323: sound1 <=  91370;
	4324: sound1 <=  119537;
	4325: sound1 <=  169373;
	4326: sound1 <=  185120;
	4327: sound1 <=  67993;
	4328: sound1 <=  53986;
	4329: sound1 <=  53894;
	4330: sound1 <=  52063;
	4331: sound1 <=  78156;
	4332: sound1 <=  136566;
	4333: sound1 <=  144775;
	4334: sound1 <=  127502;
	4335: sound1 <=  137543;
	4336: sound1 <=  131226;
	4337: sound1 <=  104279;
	4338: sound1 <=  104828;
	4339: sound1 <=  117767;
	4340: sound1 <=  94910;
	4341: sound1 <=  52368;
	4342: sound1 <=  57709;
	4343: sound1 <=  137512;
	4344: sound1 <=  174652;
	4345: sound1 <=  183075;
	4346: sound1 <=  203278;
	4347: sound1 <=  197052;
	4348: sound1 <=  186829;
	4349: sound1 <=  23621;
	4350: sound1 <=  -63354;
	4351: sound1 <=  -71564;
	4352: sound1 <=  -95398;
	4353: sound1 <=  -128998;
	4354: sound1 <=  -115967;
	4355: sound1 <=  -59662;
	4356: sound1 <=  -9186;
	4357: sound1 <=  33875;
	4358: sound1 <=  87982;
	4359: sound1 <=  161926;
	4360: sound1 <=  211670;
	4361: sound1 <=  236115;
	4362: sound1 <=  261047;
	4363: sound1 <=  135986;
	4364: sound1 <=  62225;
	4365: sound1 <=  87585;
	4366: sound1 <=  111389;
	4367: sound1 <=  143005;
	4368: sound1 <=  179932;
	4369: sound1 <=  216827;
	4370: sound1 <=  224915;
	4371: sound1 <=  247070;
	4372: sound1 <=  190491;
	4373: sound1 <=  70709;
	4374: sound1 <=  91339;
	4375: sound1 <=  84900;
	4376: sound1 <=  44830;
	4377: sound1 <=  26031;
	4378: sound1 <=  54871;
	4379: sound1 <=  101196;
	4380: sound1 <=  136871;
	4381: sound1 <=  148499;
	4382: sound1 <=  162048;
	4383: sound1 <=  157837;
	4384: sound1 <=  179077;
	4385: sound1 <=  66650;
	4386: sound1 <=  -39673;
	4387: sound1 <=  -72540;
	4388: sound1 <=  -107269;
	4389: sound1 <=  -69366;
	4390: sound1 <=  -24658;
	4391: sound1 <=  -32898;
	4392: sound1 <=  -116394;
	4393: sound1 <=  -69305;
	4394: sound1 <=  -27191;
	4395: sound1 <=  16724;
	4396: sound1 <=  50049;
	4397: sound1 <=  -49713;
	4398: sound1 <=  -102661;
	4399: sound1 <=  -119751;
	4400: sound1 <=  -71381;
	4401: sound1 <=  549;
	4402: sound1 <=  37445;
	4403: sound1 <=  73059;
	4404: sound1 <=  88867;
	4405: sound1 <=  -30060;
	4406: sound1 <=  -76233;
	4407: sound1 <=  -67505;
	4408: sound1 <=  -86426;
	4409: sound1 <=  -100098;
	4410: sound1 <=  -93048;
	4411: sound1 <=  -55481;
	4412: sound1 <=  -9369;
	4413: sound1 <=  -31;
	4414: sound1 <=  23163;
	4415: sound1 <=  67230;
	4416: sound1 <=  106384;
	4417: sound1 <=  157227;
	4418: sound1 <=  200653;
	4419: sound1 <=  216553;
	4420: sound1 <=  205841;
	4421: sound1 <=  83221;
	4422: sound1 <=  -11353;
	4423: sound1 <=  -68024;
	4424: sound1 <=  -66010;
	4425: sound1 <=  -32013;
	4426: sound1 <=  916;
	4427: sound1 <=  68695;
	4428: sound1 <=  102570;
	4429: sound1 <=  123322;
	4430: sound1 <=  90668;
	4431: sound1 <=  -64880;
	4432: sound1 <=  -87799;
	4433: sound1 <=  -81604;
	4434: sound1 <=  -55756;
	4435: sound1 <=  -16113;
	4436: sound1 <=  -11414;
	4437: sound1 <=  3632;
	4438: sound1 <=  18616;
	4439: sound1 <=  12756;
	4440: sound1 <=  7843;
	4441: sound1 <=  -2411;
	4442: sound1 <=  23926;
	4443: sound1 <=  62531;
	4444: sound1 <=  104736;
	4445: sound1 <=  16602;
	4446: sound1 <=  -58411;
	4447: sound1 <=  -28503;
	4448: sound1 <=  -336;
	4449: sound1 <=  41168;
	4450: sound1 <=  65399;
	4451: sound1 <=  78491;
	4452: sound1 <=  96771;
	4453: sound1 <=  115875;
	4454: sound1 <=  94788;
	4455: sound1 <=  104858;
	4456: sound1 <=  148651;
	4457: sound1 <=  178467;
	4458: sound1 <=  172668;
	4459: sound1 <=  181213;
	4460: sound1 <=  216675;
	4461: sound1 <=  235016;
	4462: sound1 <=  255615;
	4463: sound1 <=  216125;
	4464: sound1 <=  87097;
	4465: sound1 <=  39429;
	4466: sound1 <=  -21790;
	4467: sound1 <=  -49072;
	4468: sound1 <=  -82092;
	4469: sound1 <=  -110657;
	4470: sound1 <=  -117554;
	4471: sound1 <=  -105988;
	4472: sound1 <=  -87524;
	4473: sound1 <=  -53680;
	4474: sound1 <=  -25513;
	4475: sound1 <=  2838;
	4476: sound1 <=  56824;
	4477: sound1 <=  94574;
	4478: sound1 <=  138794;
	4479: sound1 <=  168549;
	4480: sound1 <=  52521;
	4481: sound1 <=  10651;
	4482: sound1 <=  13397;
	4483: sound1 <=  25543;
	4484: sound1 <=  33997;
	4485: sound1 <=  38177;
	4486: sound1 <=  25055;
	4487: sound1 <=  -16632;
	4488: sound1 <=  -11108;
	4489: sound1 <=  -18646;
	4490: sound1 <=  -39856;
	4491: sound1 <=  -73669;
	4492: sound1 <=  -114258;
	4493: sound1 <=  -145386;
	4494: sound1 <=  -139648;
	4495: sound1 <=  -115753;
	4496: sound1 <=  -79834;
	4497: sound1 <=  -12054;
	4498: sound1 <=  27100;
	4499: sound1 <=  32104;
	4500: sound1 <=  60852;
	4501: sound1 <=  99823;
	4502: sound1 <=  112701;
	4503: sound1 <=  116486;
	4504: sound1 <=  104248;
	4505: sound1 <=  98633;
	4506: sound1 <=  64545;
	4507: sound1 <=  -122162;
	4508: sound1 <=  -190277;
	4509: sound1 <=  -205963;
	4510: sound1 <=  -216217;
	4511: sound1 <=  -219299;
	4512: sound1 <=  -201050;
	4513: sound1 <=  -192383;
	4514: sound1 <=  -172821;
	4515: sound1 <=  -108582;
	4516: sound1 <=  -25116;
	4517: sound1 <=  17395;
	4518: sound1 <=  19928;
	4519: sound1 <=  9064;
	4520: sound1 <=  14587;
	4521: sound1 <=  7019;
	4522: sound1 <=  -12085;
	4523: sound1 <=  -28442;
	4524: sound1 <=  -46112;
	4525: sound1 <=  -15015;
	4526: sound1 <=  33997;
	4527: sound1 <=  51910;
	4528: sound1 <=  64270;
	4529: sound1 <=  28320;
	4530: sound1 <=  7233;
	4531: sound1 <=  -124695;
	4532: sound1 <=  -205963;
	4533: sound1 <=  -198395;
	4534: sound1 <=  -188873;
	4535: sound1 <=  -210754;
	4536: sound1 <=  -208038;
	4537: sound1 <=  -183716;
	4538: sound1 <=  -150574;
	4539: sound1 <=  -100189;
	4540: sound1 <=  -70526;
	4541: sound1 <=  -53589;
	4542: sound1 <=  -17365;
	4543: sound1 <=  22491;
	4544: sound1 <=  4639;
	4545: sound1 <=  -2502;
	4546: sound1 <=  10773;
	4547: sound1 <=  35248;
	4548: sound1 <=  73914;
	4549: sound1 <=  105957;
	4550: sound1 <=  118530;
	4551: sound1 <=  115967;
	4552: sound1 <=  133820;
	4553: sound1 <=  160797;
	4554: sound1 <=  181671;
	4555: sound1 <=  175507;
	4556: sound1 <=  189575;
	4557: sound1 <=  188751;
	4558: sound1 <=  217316;
	4559: sound1 <=  257263;
	4560: sound1 <=  284302;
	4561: sound1 <=  288300;
	4562: sound1 <=  238556;
	4563: sound1 <=  212067;
	4564: sound1 <=  195709;
	4565: sound1 <=  190033;
	4566: sound1 <=  192047;
	4567: sound1 <=  183380;
	4568: sound1 <=  177826;
	4569: sound1 <=  180542;
	4570: sound1 <=  164825;
	4571: sound1 <=  146088;
	4572: sound1 <=  159515;
	4573: sound1 <=  190063;
	4574: sound1 <=  197418;
	4575: sound1 <=  183289;
	4576: sound1 <=  145142;
	4577: sound1 <=  104065;
	4578: sound1 <=  67413;
	4579: sound1 <=  51666;
	4580: sound1 <=  28564;
	4581: sound1 <=  -1770;
	4582: sound1 <=  4333;
	4583: sound1 <=  71594;
	4584: sound1 <=  131500;
	4585: sound1 <=  130219;
	4586: sound1 <=  113922;
	4587: sound1 <=  88470;
	4588: sound1 <=  71930;
	4589: sound1 <=  68085;
	4590: sound1 <=  51147;
	4591: sound1 <=  10803;
	4592: sound1 <=  -23712;
	4593: sound1 <=  11322;
	4594: sound1 <=  43274;
	4595: sound1 <=  41138;
	4596: sound1 <=  -101349;
	4597: sound1 <=  -204559;
	4598: sound1 <=  -251282;
	4599: sound1 <=  -326874;
	4600: sound1 <=  -310669;
	4601: sound1 <=  -303467;
	4602: sound1 <=  -283051;
	4603: sound1 <=  -236847;
	4604: sound1 <=  -185303;
	4605: sound1 <=  -123474;
	4606: sound1 <=  -72998;
	4607: sound1 <=  -32104;
	4608: sound1 <=  15594;
	4609: sound1 <=  -9613;
	4610: sound1 <=  70099;
	4611: sound1 <=  131836;
	4612: sound1 <=  125458;
	4613: sound1 <=  32288;
	4614: sound1 <=  79712;
	4615: sound1 <=  130615;
	4616: sound1 <=  196930;
	4617: sound1 <=  193939;
	4618: sound1 <=  88684;
	4619: sound1 <=  74158;
	4620: sound1 <=  52246;
	4621: sound1 <=  43091;
	4622: sound1 <=  31067;
	4623: sound1 <=  40283;
	4624: sound1 <=  50049;
	4625: sound1 <=  59723;
	4626: sound1 <=  29510;
	4627: sound1 <=  -7751;
	4628: sound1 <=  37109;
	4629: sound1 <=  63446;
	4630: sound1 <=  81970;
	4631: sound1 <=  33203;
	4632: sound1 <=  -95642;
	4633: sound1 <=  -87677;
	4634: sound1 <=  -101135;
	4635: sound1 <=  -120178;
	4636: sound1 <=  -126190;
	4637: sound1 <=  -151672;
	4638: sound1 <=  -134155;
	4639: sound1 <=  -122528;
	4640: sound1 <=  -99670;
	4641: sound1 <=  -56030;
	4642: sound1 <=  -17731;
	4643: sound1 <=  45380;
	4644: sound1 <=  99670;
	4645: sound1 <=  112671;
	4646: sound1 <=  145172;
	4647: sound1 <=  191833;
	4648: sound1 <=  234985;
	4649: sound1 <=  262451;
	4650: sound1 <=  155060;
	4651: sound1 <=  116730;
	4652: sound1 <=  87524;
	4653: sound1 <=  80292;
	4654: sound1 <=  97809;
	4655: sound1 <=  115662;
	4656: sound1 <=  158203;
	4657: sound1 <=  182861;
	4658: sound1 <=  196228;
	4659: sound1 <=  234070;
	4660: sound1 <=  206635;
	4661: sound1 <=  86151;
	4662: sound1 <=  78491;
	4663: sound1 <=  84869;
	4664: sound1 <=  118317;
	4665: sound1 <=  139099;
	4666: sound1 <=  161774;
	4667: sound1 <=  195557;
	4668: sound1 <=  202240;
	4669: sound1 <=  200592;
	4670: sound1 <=  199982;
	4671: sound1 <=  130066;
	4672: sound1 <=  -96802;
	4673: sound1 <=  -138245;
	4674: sound1 <=  -173370;
	4675: sound1 <=  -201782;
	4676: sound1 <=  -215942;
	4677: sound1 <=  -217804;
	4678: sound1 <=  -206482;
	4679: sound1 <=  -190033;
	4680: sound1 <=  -162872;
	4681: sound1 <=  -153809;
	4682: sound1 <=  -142120;
	4683: sound1 <=  -80811;
	4684: sound1 <=  -15411;
	4685: sound1 <=  10529;
	4686: sound1 <=  52368;
	4687: sound1 <=  64484;
	4688: sound1 <=  104736;
	4689: sound1 <=  130066;
	4690: sound1 <=  152191;
	4691: sound1 <=  190521;
	4692: sound1 <=  177551;
	4693: sound1 <=  166351;
	4694: sound1 <=  155579;
	4695: sound1 <=  126099;
	4696: sound1 <=  89081;
	4697: sound1 <=  77606;
	4698: sound1 <=  100067;
	4699: sound1 <=  146301;
	4700: sound1 <=  211975;
	4701: sound1 <=  290161;
	4702: sound1 <=  316193;
	4703: sound1 <=  326019;
	4704: sound1 <=  312408;
	4705: sound1 <=  277222;
	4706: sound1 <=  274384;
	4707: sound1 <=  269318;
	4708: sound1 <=  265320;
	4709: sound1 <=  270203;
	4710: sound1 <=  257050;
	4711: sound1 <=  223602;
	4712: sound1 <=  203827;
	4713: sound1 <=  195068;
	4714: sound1 <=  187531;
	4715: sound1 <=  171997;
	4716: sound1 <=  147949;
	4717: sound1 <=  97504;
	4718: sound1 <=  71381;
	4719: sound1 <=  70129;
	4720: sound1 <=  33234;
	4721: sound1 <=  -23407;
	4722: sound1 <=  -60028;
	4723: sound1 <=  -55389;
	4724: sound1 <=  -89203;
	4725: sound1 <=  -129395;
	4726: sound1 <=  -141602;
	4727: sound1 <=  -150513;
	4728: sound1 <=  -171539;
	4729: sound1 <=  -200409;
	4730: sound1 <=  -241547;
	4731: sound1 <=  -270447;
	4732: sound1 <=  -238983;
	4733: sound1 <=  -197662;
	4734: sound1 <=  -159332;
	4735: sound1 <=  -161041;
	4736: sound1 <=  -151337;
	4737: sound1 <=  -163818;
	4738: sound1 <=  -165192;
	4739: sound1 <=  -129181;
	4740: sound1 <=  -108643;
	4741: sound1 <=  -85236;
	4742: sound1 <=  -32867;
	4743: sound1 <=  -24017;
	4744: sound1 <=  -54047;
	4745: sound1 <=  -67200;
	4746: sound1 <=  -65491;
	4747: sound1 <=  -75317;
	4748: sound1 <=  -80139;
	4749: sound1 <=  -82214;
	4750: sound1 <=  -89081;
	4751: sound1 <=  -81940;
	4752: sound1 <=  -69031;
	4753: sound1 <=  -84991;
	4754: sound1 <=  -76050;
	4755: sound1 <=  -66467;
	4756: sound1 <=  -80994;
	4757: sound1 <=  -85693;
	4758: sound1 <=  -71747;
	4759: sound1 <=  -75073;
	4760: sound1 <=  -106995;
	4761: sound1 <=  -84991;
	4762: sound1 <=  -89203;
	4763: sound1 <=  -109009;
	4764: sound1 <=  -93292;
	4765: sound1 <=  -56030;
	4766: sound1 <=  -26093;
	4767: sound1 <=  -5707;
	4768: sound1 <=  -55817;
	4769: sound1 <=  -171448;
	4770: sound1 <=  -174957;
	4771: sound1 <=  -176239;
	4772: sound1 <=  -182343;
	4773: sound1 <=  -187561;
	4774: sound1 <=  -176300;
	4775: sound1 <=  -155548;
	4776: sound1 <=  -91003;
	4777: sound1 <=  -23926;
	4778: sound1 <=  8911;
	4779: sound1 <=  12665;
	4780: sound1 <=  20782;
	4781: sound1 <=  50629;
	4782: sound1 <=  53711;
	4783: sound1 <=  64880;
	4784: sound1 <=  93719;
	4785: sound1 <=  120209;
	4786: sound1 <=  118896;
	4787: sound1 <=  138489;
	4788: sound1 <=  158661;
	4789: sound1 <=  76324;
	4790: sound1 <=  99121;
	4791: sound1 <=  140808;
	4792: sound1 <=  173523;
	4793: sound1 <=  230225;
	4794: sound1 <=  264374;
	4795: sound1 <=  262787;
	4796: sound1 <=  226440;
	4797: sound1 <=  209106;
	4798: sound1 <=  188843;
	4799: sound1 <=  219727;
	4800: sound1 <=  127014;
	4801: sound1 <=  21912;
	4802: sound1 <=  -3296;
	4803: sound1 <=  -38666;
	4804: sound1 <=  -34729;
	4805: sound1 <=  -24994;
	4806: sound1 <=  -43152;
	4807: sound1 <=  -49774;
	4808: sound1 <=  -55908;
	4809: sound1 <=  -45868;
	4810: sound1 <=  -38025;
	4811: sound1 <=  -46722;
	4812: sound1 <=  -60028;
	4813: sound1 <=  -37720;
	4814: sound1 <=  7690;
	4815: sound1 <=  69336;
	4816: sound1 <=  114197;
	4817: sound1 <=  130035;
	4818: sound1 <=  135071;
	4819: sound1 <=  153870;
	4820: sound1 <=  196167;
	4821: sound1 <=  167908;
	4822: sound1 <=  28351;
	4823: sound1 <=  -4944;
	4824: sound1 <=  -11536;
	4825: sound1 <=  -14130;
	4826: sound1 <=  6256;
	4827: sound1 <=  48981;
	4828: sound1 <=  79529;
	4829: sound1 <=  152496;
	4830: sound1 <=  206665;
	4831: sound1 <=  242065;
	4832: sound1 <=  258850;
	4833: sound1 <=  277649;
	4834: sound1 <=  144165;
	4835: sound1 <=  13184;
	4836: sound1 <=  -8636;
	4837: sound1 <=  -67810;
	4838: sound1 <=  -75012;
	4839: sound1 <=  -102875;
	4840: sound1 <=  -111572;
	4841: sound1 <=  -80688;
	4842: sound1 <=  -28229;
	4843: sound1 <=  -1556;
	4844: sound1 <=  -1526;
	4845: sound1 <=  -1495;
	4846: sound1 <=  28992;
	4847: sound1 <=  81726;
	4848: sound1 <=  138123;
	4849: sound1 <=  182617;
	4850: sound1 <=  212463;
	4851: sound1 <=  277924;
	4852: sound1 <=  331451;
	4853: sound1 <=  329651;
	4854: sound1 <=  329987;
	4855: sound1 <=  352631;
	4856: sound1 <=  364441;
	4857: sound1 <=  341034;
	4858: sound1 <=  331207;
	4859: sound1 <=  339264;
	4860: sound1 <=  355530;
	4861: sound1 <=  340332;
	4862: sound1 <=  314392;
	4863: sound1 <=  310516;
	4864: sound1 <=  293640;
	4865: sound1 <=  243347;
	4866: sound1 <=  224884;
	4867: sound1 <=  240204;
	4868: sound1 <=  229218;
	4869: sound1 <=  214417;
	4870: sound1 <=  207001;
	4871: sound1 <=  175568;
	4872: sound1 <=  155914;
	4873: sound1 <=  92682;
	4874: sound1 <=  -67505;
	4875: sound1 <=  -112549;
	4876: sound1 <=  -167816;
	4877: sound1 <=  -203583;
	4878: sound1 <=  -268341;
	4879: sound1 <=  -345398;
	4880: sound1 <=  -391876;
	4881: sound1 <=  -408569;
	4882: sound1 <=  -409821;
	4883: sound1 <=  -396729;
	4884: sound1 <=  -332031;
	4885: sound1 <=  -283630;
	4886: sound1 <=  -227295;
	4887: sound1 <=  -163025;
	4888: sound1 <=  -120850;
	4889: sound1 <=  -104187;
	4890: sound1 <=  -63049;
	4891: sound1 <=  -15533;
	4892: sound1 <=  -129181;
	4893: sound1 <=  -186401;
	4894: sound1 <=  -156830;
	4895: sound1 <=  -153107;
	4896: sound1 <=  -163177;
	4897: sound1 <=  -132019;
	4898: sound1 <=  -88196;
	4899: sound1 <=  -14679;
	4900: sound1 <=  50415;
	4901: sound1 <=  -5402;
	4902: sound1 <=  -102600;
	4903: sound1 <=  -102325;
	4904: sound1 <=  -126892;
	4905: sound1 <=  -126282;
	4906: sound1 <=  -127991;
	4907: sound1 <=  -129822;
	4908: sound1 <=  -156128;
	4909: sound1 <=  -247162;
	4910: sound1 <=  -199371;
	4911: sound1 <=  -144562;
	4912: sound1 <=  -108307;
	4913: sound1 <=  -62897;
	4914: sound1 <=  -21545;
	4915: sound1 <=  -93811;
	4916: sound1 <=  -118439;
	4917: sound1 <=  -76324;
	4918: sound1 <=  -19226;
	4919: sound1 <=  31677;
	4920: sound1 <=  86090;
	4921: sound1 <=  18036;
	4922: sound1 <=  -15991;
	4923: sound1 <=  45624;
	4924: sound1 <=  132568;
	4925: sound1 <=  208984;
	4926: sound1 <=  228485;
	4927: sound1 <=  258240;
	4928: sound1 <=  125946;
	4929: sound1 <=  122406;
	4930: sound1 <=  161957;
	4931: sound1 <=  203064;
	4932: sound1 <=  155426;
	4933: sound1 <=  169098;
	4934: sound1 <=  203613;
	4935: sound1 <=  172394;
	4936: sound1 <=  89020;
	4937: sound1 <=  145966;
	4938: sound1 <=  149323;
	4939: sound1 <=  167297;
	4940: sound1 <=  212158;
	4941: sound1 <=  237701;
	4942: sound1 <=  139923;
	4943: sound1 <=  154694;
	4944: sound1 <=  241211;
	4945: sound1 <=  254395;
	4946: sound1 <=  274200;
	4947: sound1 <=  139435;
	4948: sound1 <=  117828;
	4949: sound1 <=  114410;
	4950: sound1 <=  56274;
	4951: sound1 <=  6378;
	4952: sound1 <=  -14404;
	4953: sound1 <=  16418;
	4954: sound1 <=  20386;
	4955: sound1 <=  35828;
	4956: sound1 <=  21576;
	4957: sound1 <=  27161;
	4958: sound1 <=  61157;
	4959: sound1 <=  84106;
	4960: sound1 <=  89600;
	4961: sound1 <=  55176;
	4962: sound1 <=  1495;
	4963: sound1 <=  -9918;
	4964: sound1 <=  12604;
	4965: sound1 <=  46143;
	4966: sound1 <=  60760;
	4967: sound1 <=  82520;
	4968: sound1 <=  65704;
	4969: sound1 <=  63416;
	4970: sound1 <=  -6775;
	4971: sound1 <=  -213776;
	4972: sound1 <=  -242249;
	4973: sound1 <=  -254059;
	4974: sound1 <=  -250671;
	4975: sound1 <=  -253357;
	4976: sound1 <=  -229797;
	4977: sound1 <=  -180328;
	4978: sound1 <=  -176605;
	4979: sound1 <=  -169067;
	4980: sound1 <=  -126190;
	4981: sound1 <=  -79834;
	4982: sound1 <=  -48340;
	4983: sound1 <=  22369;
	4984: sound1 <=  97748;
	4985: sound1 <=  154694;
	4986: sound1 <=  193298;
	4987: sound1 <=  237640;
	4988: sound1 <=  291687;
	4989: sound1 <=  292755;
	4990: sound1 <=  326721;
	4991: sound1 <=  338379;
	4992: sound1 <=  338593;
	4993: sound1 <=  348511;
	4994: sound1 <=  372772;
	4995: sound1 <=  363007;
	4996: sound1 <=  356720;
	4997: sound1 <=  285767;
	4998: sound1 <=  173767;
	4999: sound1 <=  172424;
	5000: sound1 <=  122223;
	5001: sound1 <=  89661;
	5002: sound1 <=  55969;
	5003: sound1 <=  39612;
	5004: sound1 <=  42328;
	5005: sound1 <=  40222;
	5006: sound1 <=  27863;
	5007: sound1 <=  28839;
	5008: sound1 <=  39124;
	5009: sound1 <=  15778;
	5010: sound1 <=  -32227;
	5011: sound1 <=  -82794;
	5012: sound1 <=  -84900;
	5013: sound1 <=  -85022;
	5014: sound1 <=  -117035;
	5015: sound1 <=  -105347;
	5016: sound1 <=  -75958;
	5017: sound1 <=  -29358;
	5018: sound1 <=  26093;
	5019: sound1 <=  43976;
	5020: sound1 <=  46265;
	5021: sound1 <=  28137;
	5022: sound1 <=  76782;
	5023: sound1 <=  119507;
	5024: sound1 <=  129486;
	5025: sound1 <=  125153;
	5026: sound1 <=  82031;
	5027: sound1 <=  100281;
	5028: sound1 <=  125305;
	5029: sound1 <=  129852;
	5030: sound1 <=  132782;
	5031: sound1 <=  118683;
	5032: sound1 <=  122040;
	5033: sound1 <=  122498;
	5034: sound1 <=  107574;
	5035: sound1 <=  93811;
	5036: sound1 <=  53864;
	5037: sound1 <=  10162;
	5038: sound1 <=  -12695;
	5039: sound1 <=  -42999;
	5040: sound1 <=  -85052;
	5041: sound1 <=  -130585;
	5042: sound1 <=  -150574;
	5043: sound1 <=  -168274;
	5044: sound1 <=  -190277;
	5045: sound1 <=  -214905;
	5046: sound1 <=  -250031;
	5047: sound1 <=  -258820;
	5048: sound1 <=  -259521;
	5049: sound1 <=  -241638;
	5050: sound1 <=  -210052;
	5051: sound1 <=  -174408;
	5052: sound1 <=  -154266;
	5053: sound1 <=  -147491;
	5054: sound1 <=  -93414;
	5055: sound1 <=  -48615;
	5056: sound1 <=  -30701;
	5057: sound1 <=  -27496;
	5058: sound1 <=  -40863;
	5059: sound1 <=  -26733;
	5060: sound1 <=  -25787;
	5061: sound1 <=  -44037;
	5062: sound1 <=  -69885;
	5063: sound1 <=  -81482;
	5064: sound1 <=  -70221;
	5065: sound1 <=  -71381;
	5066: sound1 <=  -99518;
	5067: sound1 <=  -99121;
	5068: sound1 <=  -112579;
	5069: sound1 <=  -147949;
	5070: sound1 <=  -164063;
	5071: sound1 <=  -158905;
	5072: sound1 <=  -158020;
	5073: sound1 <=  -192444;
	5074: sound1 <=  -229370;
	5075: sound1 <=  -207520;
	5076: sound1 <=  -194061;
	5077: sound1 <=  -157166;
	5078: sound1 <=  -120911;
	5079: sound1 <=  -109283;
	5080: sound1 <=  -102020;
	5081: sound1 <=  -87463;
	5082: sound1 <=  -39215;
	5083: sound1 <=  20020;
	5084: sound1 <=  37048;
	5085: sound1 <=  60760;
	5086: sound1 <=  65216;
	5087: sound1 <=  102448;
	5088: sound1 <=  126282;
	5089: sound1 <=  91003;
	5090: sound1 <=  108643;
	5091: sound1 <=  158569;
	5092: sound1 <=  192657;
	5093: sound1 <=  247009;
	5094: sound1 <=  257813;
	5095: sound1 <=  254211;
	5096: sound1 <=  215393;
	5097: sound1 <=  215881;
	5098: sound1 <=  233307;
	5099: sound1 <=  193817;
	5100: sound1 <=  176392;
	5101: sound1 <=  176270;
	5102: sound1 <=  154968;
	5103: sound1 <=  155243;
	5104: sound1 <=  170868;
	5105: sound1 <=  174194;
	5106: sound1 <=  174316;
	5107: sound1 <=  175476;
	5108: sound1 <=  202484;
	5109: sound1 <=  217377;
	5110: sound1 <=  219482;
	5111: sound1 <=  195801;
	5112: sound1 <=  177368;
	5113: sound1 <=  184418;
	5114: sound1 <=  207428;
	5115: sound1 <=  221100;
	5116: sound1 <=  221008;
	5117: sound1 <=  218719;
	5118: sound1 <=  232056;
	5119: sound1 <=  245941;
	5120: sound1 <=  225769;
	5121: sound1 <=  161072;
	5122: sound1 <=  135071;
	5123: sound1 <=  139038;
	5124: sound1 <=  123840;
	5125: sound1 <=  101288;
	5126: sound1 <=  60669;
	5127: sound1 <=  31342;
	5128: sound1 <=  -2197;
	5129: sound1 <=  -27222;
	5130: sound1 <=  -27924;
	5131: sound1 <=  -15717;
	5132: sound1 <=  -36591;
	5133: sound1 <=  -75012;
	5134: sound1 <=  -64850;
	5135: sound1 <=  -29694;
	5136: sound1 <=  -24536;
	5137: sound1 <=  -17334;
	5138: sound1 <=  -7843;
	5139: sound1 <=  -22491;
	5140: sound1 <=  -4578;
	5141: sound1 <=  8606;
	5142: sound1 <=  -4974;
	5143: sound1 <=  -28687;
	5144: sound1 <=  -49561;
	5145: sound1 <=  -42206;
	5146: sound1 <=  -21423;
	5147: sound1 <=  11536;
	5148: sound1 <=  48309;
	5149: sound1 <=  82001;
	5150: sound1 <=  80353;
	5151: sound1 <=  62408;
	5152: sound1 <=  41077;
	5153: sound1 <=  40436;
	5154: sound1 <=  61890;
	5155: sound1 <=  66895;
	5156: sound1 <=  52002;
	5157: sound1 <=  31952;
	5158: sound1 <=  64392;
	5159: sound1 <=  73822;
	5160: sound1 <=  66284;
	5161: sound1 <=  37018;
	5162: sound1 <=  -12573;
	5163: sound1 <=  -27069;
	5164: sound1 <=  -18219;
	5165: sound1 <=  -28076;
	5166: sound1 <=  -37048;
	5167: sound1 <=  -67993;
	5168: sound1 <=  -72357;
	5169: sound1 <=  -86670;
	5170: sound1 <=  -76172;
	5171: sound1 <=  -47882;
	5172: sound1 <=  -27100;
	5173: sound1 <=  -13397;
	5174: sound1 <=  3265;
	5175: sound1 <=  4059;
	5176: sound1 <=  17426;
	5177: sound1 <=  19775;
	5178: sound1 <=  20538;
	5179: sound1 <=  53253;
	5180: sound1 <=  89966;
	5181: sound1 <=  115631;
	5182: sound1 <=  144928;
	5183: sound1 <=  159393;
	5184: sound1 <=  163330;
	5185: sound1 <=  137909;
	5186: sound1 <=  136719;
	5187: sound1 <=  59143;
	5188: sound1 <=  -100525;
	5189: sound1 <=  -115906;
	5190: sound1 <=  -116638;
	5191: sound1 <=  -148926;
	5192: sound1 <=  -188965;
	5193: sound1 <=  -223785;
	5194: sound1 <=  -225983;
	5195: sound1 <=  -218506;
	5196: sound1 <=  -216766;
	5197: sound1 <=  -228302;
	5198: sound1 <=  -218079;
	5199: sound1 <=  -180328;
	5200: sound1 <=  -129456;
	5201: sound1 <=  -98419;
	5202: sound1 <=  -65643;
	5203: sound1 <=  -12939;
	5204: sound1 <=  51331;
	5205: sound1 <=  98602;
	5206: sound1 <=  166107;
	5207: sound1 <=  211761;
	5208: sound1 <=  203766;
	5209: sound1 <=  192505;
	5210: sound1 <=  205933;
	5211: sound1 <=  226196;
	5212: sound1 <=  239685;
	5213: sound1 <=  285156;
	5214: sound1 <=  332794;
	5215: sound1 <=  329834;
	5216: sound1 <=  306946;
	5217: sound1 <=  269379;
	5218: sound1 <=  248413;
	5219: sound1 <=  238129;
	5220: sound1 <=  234741;
	5221: sound1 <=  226868;
	5222: sound1 <=  224915;
	5223: sound1 <=  221863;
	5224: sound1 <=  227600;
	5225: sound1 <=  198334;
	5226: sound1 <=  192139;
	5227: sound1 <=  204895;
	5228: sound1 <=  197235;
	5229: sound1 <=  176178;
	5230: sound1 <=  153473;
	5231: sound1 <=  115173;
	5232: sound1 <=  91827;
	5233: sound1 <=  85022;
	5234: sound1 <=  67169;
	5235: sound1 <=  69427;
	5236: sound1 <=  88776;
	5237: sound1 <=  69397;
	5238: sound1 <=  -6287;
	5239: sound1 <=  -66528;
	5240: sound1 <=  -113708;
	5241: sound1 <=  -163910;
	5242: sound1 <=  -170898;
	5243: sound1 <=  -154602;
	5244: sound1 <=  -130768;
	5245: sound1 <=  -111603;
	5246: sound1 <=  -87189;
	5247: sound1 <=  -95215;
	5248: sound1 <=  -99060;
	5249: sound1 <=  -80536;
	5250: sound1 <=  -86212;
	5251: sound1 <=  -76660;
	5252: sound1 <=  -80658;
	5253: sound1 <=  -90729;
	5254: sound1 <=  -113373;
	5255: sound1 <=  -124786;
	5256: sound1 <=  -111816;
	5257: sound1 <=  -123413;
	5258: sound1 <=  -154358;
	5259: sound1 <=  -157471;
	5260: sound1 <=  -175812;
	5261: sound1 <=  -193512;
	5262: sound1 <=  -170441;
	5263: sound1 <=  -134094;
	5264: sound1 <=  -125580;
	5265: sound1 <=  -118591;
	5266: sound1 <=  -161926;
	5267: sound1 <=  -235443;
	5268: sound1 <=  -242401;
	5269: sound1 <=  -251556;
	5270: sound1 <=  -285950;
	5271: sound1 <=  -290039;
	5272: sound1 <=  -290009;
	5273: sound1 <=  -269012;
	5274: sound1 <=  -243042;
	5275: sound1 <=  -226776;
	5276: sound1 <=  -203552;
	5277: sound1 <=  -216339;
	5278: sound1 <=  -233765;
	5279: sound1 <=  -226868;
	5280: sound1 <=  -195496;
	5281: sound1 <=  -140137;
	5282: sound1 <=  -60150;
	5283: sound1 <=  14709;
	5284: sound1 <=  79102;
	5285: sound1 <=  147461;
	5286: sound1 <=  203918;
	5287: sound1 <=  238403;
	5288: sound1 <=  261261;
	5289: sound1 <=  156403;
	5290: sound1 <=  84930;
	5291: sound1 <=  66986;
	5292: sound1 <=  68542;
	5293: sound1 <=  89752;
	5294: sound1 <=  139923;
	5295: sound1 <=  202728;
	5296: sound1 <=  211426;
	5297: sound1 <=  198120;
	5298: sound1 <=  212128;
	5299: sound1 <=  248566;
	5300: sound1 <=  162109;
	5301: sound1 <=  115997;
	5302: sound1 <=  137085;
	5303: sound1 <=  124481;
	5304: sound1 <=  147644;
	5305: sound1 <=  69336;
	5306: sound1 <=  30151;
	5307: sound1 <=  74524;
	5308: sound1 <=  126068;
	5309: sound1 <=  159851;
	5310: sound1 <=  177734;
	5311: sound1 <=  107422;
	5312: sound1 <=  127655;
	5313: sound1 <=  230408;
	5314: sound1 <=  219666;
	5315: sound1 <=  187378;
	5316: sound1 <=  245667;
	5317: sound1 <=  294189;
	5318: sound1 <=  315796;
	5319: sound1 <=  270721;
	5320: sound1 <=  122589;
	5321: sound1 <=  89203;
	5322: sound1 <=  62439;
	5323: sound1 <=  54749;
	5324: sound1 <=  56702;
	5325: sound1 <=  36316;
	5326: sound1 <=  40924;
	5327: sound1 <=  41779;
	5328: sound1 <=  67352;
	5329: sound1 <=  115234;
	5330: sound1 <=  69153;
	5331: sound1 <=  55084;
	5332: sound1 <=  16357;
	5333: sound1 <=  -60059;
	5334: sound1 <=  -19135;
	5335: sound1 <=  -9003;
	5336: sound1 <=  11841;
	5337: sound1 <=  63965;
	5338: sound1 <=  106506;
	5339: sound1 <=  159882;
	5340: sound1 <=  97107;
	5341: sound1 <=  67596;
	5342: sound1 <=  86945;
	5343: sound1 <=  54871;
	5344: sound1 <=  35034;
	5345: sound1 <=  22278;
	5346: sound1 <=  23010;
	5347: sound1 <=  28839;
	5348: sound1 <=  41687;
	5349: sound1 <=  53833;
	5350: sound1 <=  66772;
	5351: sound1 <=  104004;
	5352: sound1 <=  159790;
	5353: sound1 <=  201843;
	5354: sound1 <=  209625;
	5355: sound1 <=  195496;
	5356: sound1 <=  161743;
	5357: sound1 <=  188507;
	5358: sound1 <=  207428;
	5359: sound1 <=  214172;
	5360: sound1 <=  250336;
	5361: sound1 <=  254303;
	5362: sound1 <=  119324;
	5363: sound1 <=  16846;
	5364: sound1 <=  -25360;
	5365: sound1 <=  -45715;
	5366: sound1 <=  14618;
	5367: sound1 <=  9308;
	5368: sound1 <=  -79987;
	5369: sound1 <=  -36713;
	5370: sound1 <=  -90942;
	5371: sound1 <=  -64117;
	5372: sound1 <=  18066;
	5373: sound1 <=  -13336;
	5374: sound1 <=  -77148;
	5375: sound1 <=  -30334;
	5376: sound1 <=  -55359;
	5377: sound1 <=  -54291;
	5378: sound1 <=  -73151;
	5379: sound1 <=  -101563;
	5380: sound1 <=  -115204;
	5381: sound1 <=  -124664;
	5382: sound1 <=  -116669;
	5383: sound1 <=  -134644;
	5384: sound1 <=  -125336;
	5385: sound1 <=  -121216;
	5386: sound1 <=  -123718;
	5387: sound1 <=  -139740;
	5388: sound1 <=  -160614;
	5389: sound1 <=  -187531;
	5390: sound1 <=  -250031;
	5391: sound1 <=  -291199;
	5392: sound1 <=  -271271;
	5393: sound1 <=  -255676;
	5394: sound1 <=  -212921;
	5395: sound1 <=  -207245;
	5396: sound1 <=  -169556;
	5397: sound1 <=  -222198;
	5398: sound1 <=  -163666;
	5399: sound1 <=  -154297;
	5400: sound1 <=  -164429;
	5401: sound1 <=  -138733;
	5402: sound1 <=  -140503;
	5403: sound1 <=  -111176;
	5404: sound1 <=  -160583;
	5405: sound1 <=  -159973;
	5406: sound1 <=  -106873;
	5407: sound1 <=  -39764;
	5408: sound1 <=  -75348;
	5409: sound1 <=  -91125;
	5410: sound1 <=  -4395;
	5411: sound1 <=  -671;
	5412: sound1 <=  77118;
	5413: sound1 <=  138611;
	5414: sound1 <=  236511;
	5415: sound1 <=  298157;
	5416: sound1 <=  273773;
	5417: sound1 <=  270691;
	5418: sound1 <=  241943;
	5419: sound1 <=  243103;
	5420: sound1 <=  220917;
	5421: sound1 <=  189178;
	5422: sound1 <=  177856;
	5423: sound1 <=  147888;
	5424: sound1 <=  164917;
	5425: sound1 <=  199951;
	5426: sound1 <=  237427;
	5427: sound1 <=  166443;
	5428: sound1 <=  147614;
	5429: sound1 <=  163696;
	5430: sound1 <=  150269;
	5431: sound1 <=  65887;
	5432: sound1 <=  21362;
	5433: sound1 <=  13153;
	5434: sound1 <=  10559;
	5435: sound1 <=  63232;
	5436: sound1 <=  24353;
	5437: sound1 <=  -51331;
	5438: sound1 <=  20294;
	5439: sound1 <=  34149;
	5440: sound1 <=  85999;
	5441: sound1 <=  120636;
	5442: sound1 <=  143616;
	5443: sound1 <=  96832;
	5444: sound1 <=  25269;
	5445: sound1 <=  56244;
	5446: sound1 <=  103607;
	5447: sound1 <=  164276;
	5448: sound1 <=  186340;
	5449: sound1 <=  82245;
	5450: sound1 <=  20111;
	5451: sound1 <=  11353;
	5452: sound1 <=  44250;
	5453: sound1 <=  108490;
	5454: sound1 <=  161499;
	5455: sound1 <=  184937;
	5456: sound1 <=  207977;
	5457: sound1 <=  83160;
	5458: sound1 <=  40375;
	5459: sound1 <=  81299;
	5460: sound1 <=  93719;
	5461: sound1 <=  66895;
	5462: sound1 <=  46356;
	5463: sound1 <=  49042;
	5464: sound1 <=  37079;
	5465: sound1 <=  47516;
	5466: sound1 <=  60211;
	5467: sound1 <=  96680;
	5468: sound1 <=  98938;
	5469: sound1 <=  103394;
	5470: sound1 <=  124084;
	5471: sound1 <=  144043;
	5472: sound1 <=  157013;
	5473: sound1 <=  173584;
	5474: sound1 <=  189301;
	5475: sound1 <=  193787;
	5476: sound1 <=  187469;
	5477: sound1 <=  178864;
	5478: sound1 <=  165436;
	5479: sound1 <=  148926;
	5480: sound1 <=  118896;
	5481: sound1 <=  97321;
	5482: sound1 <=  94696;
	5483: sound1 <=  142426;
	5484: sound1 <=  151703;
	5485: sound1 <=  152374;
	5486: sound1 <=  148773;
	5487: sound1 <=  116943;
	5488: sound1 <=  99152;
	5489: sound1 <=  115967;
	5490: sound1 <=  124146;
	5491: sound1 <=  112213;
	5492: sound1 <=  -35217;
	5493: sound1 <=  -143280;
	5494: sound1 <=  -168762;
	5495: sound1 <=  -188812;
	5496: sound1 <=  -202759;
	5497: sound1 <=  -222961;
	5498: sound1 <=  -217804;
	5499: sound1 <=  -222595;
	5500: sound1 <=  -210876;
	5501: sound1 <=  -182465;
	5502: sound1 <=  -156464;
	5503: sound1 <=  -148621;
	5504: sound1 <=  -136932;
	5505: sound1 <=  -124176;
	5506: sound1 <=  -136047;
	5507: sound1 <=  -165955;
	5508: sound1 <=  -161407;
	5509: sound1 <=  -85938;
	5510: sound1 <=  -18066;
	5511: sound1 <=  29480;
	5512: sound1 <=  61676;
	5513: sound1 <=  63934;
	5514: sound1 <=  52032;
	5515: sound1 <=  70709;
	5516: sound1 <=  96436;
	5517: sound1 <=  131744;
	5518: sound1 <=  132629;
	5519: sound1 <=  112183;
	5520: sound1 <=  118958;
	5521: sound1 <=  114655;
	5522: sound1 <=  99548;
	5523: sound1 <=  104675;
	5524: sound1 <=  97717;
	5525: sound1 <=  57526;
	5526: sound1 <=  -5188;
	5527: sound1 <=  -35065;
	5528: sound1 <=  -73853;
	5529: sound1 <=  -105103;
	5530: sound1 <=  -95367;
	5531: sound1 <=  -84595;
	5532: sound1 <=  -62073;
	5533: sound1 <=  -20782;
	5534: sound1 <=  4761;
	5535: sound1 <=  7965;
	5536: sound1 <=  -37048;
	5537: sound1 <=  -49103;
	5538: sound1 <=  -56610;
	5539: sound1 <=  -65460;
	5540: sound1 <=  -74005;
	5541: sound1 <=  -78613;
	5542: sound1 <=  -74432;
	5543: sound1 <=  -36957;
	5544: sound1 <=  26306;
	5545: sound1 <=  51636;
	5546: sound1 <=  42877;
	5547: sound1 <=  36407;
	5548: sound1 <=  30029;
	5549: sound1 <=  27374;
	5550: sound1 <=  3143;
	5551: sound1 <=  -14160;
	5552: sound1 <=  -31525;
	5553: sound1 <=  -36804;
	5554: sound1 <=  -1740;
	5555: sound1 <=  15686;
	5556: sound1 <=  916;
	5557: sound1 <=  42664;
	5558: sound1 <=  97626;
	5559: sound1 <=  103058;
	5560: sound1 <=  72784;
	5561: sound1 <=  21454;
	5562: sound1 <=  13062;
	5563: sound1 <=  -8362;
	5564: sound1 <=  -8484;
	5565: sound1 <=  519;
	5566: sound1 <=  14160;
	5567: sound1 <=  10193;
	5568: sound1 <=  3357;
	5569: sound1 <=  47211;
	5570: sound1 <=  83710;
	5571: sound1 <=  79254;
	5572: sound1 <=  65491;
	5573: sound1 <=  63873;
	5574: sound1 <=  43030;
	5575: sound1 <=  19928;
	5576: sound1 <=  -12756;
	5577: sound1 <=  -21027;
	5578: sound1 <=  -25482;
	5579: sound1 <=  -31921;
	5580: sound1 <=  -26855;
	5581: sound1 <=  -61554;
	5582: sound1 <=  -97473;
	5583: sound1 <=  -90302;
	5584: sound1 <=  -120361;
	5585: sound1 <=  -174377;
	5586: sound1 <=  -193512;
	5587: sound1 <=  -203125;
	5588: sound1 <=  -229553;
	5589: sound1 <=  -251129;
	5590: sound1 <=  -228973;
	5591: sound1 <=  -229248;
	5592: sound1 <=  -212402;
	5593: sound1 <=  -197235;
	5594: sound1 <=  -186249;
	5595: sound1 <=  -144012;
	5596: sound1 <=  -77911;
	5597: sound1 <=  671;
	5598: sound1 <=  90881;
	5599: sound1 <=  187958;
	5600: sound1 <=  244812;
	5601: sound1 <=  299683;
	5602: sound1 <=  360687;
	5603: sound1 <=  409027;
	5604: sound1 <=  432709;
	5605: sound1 <=  458099;
	5606: sound1 <=  488953;
	5607: sound1 <=  514618;
	5608: sound1 <=  516357;
	5609: sound1 <=  483643;
	5610: sound1 <=  462555;
	5611: sound1 <=  411896;
	5612: sound1 <=  395111;
	5613: sound1 <=  364746;
	5614: sound1 <=  328796;
	5615: sound1 <=  189178;
	5616: sound1 <=  16235;
	5617: sound1 <=  -32013;
	5618: sound1 <=  -133942;
	5619: sound1 <=  -199402;
	5620: sound1 <=  -216644;
	5621: sound1 <=  -228760;
	5622: sound1 <=  -210999;
	5623: sound1 <=  -137054;
	5624: sound1 <=  -104126;
	5625: sound1 <=  -95337;
	5626: sound1 <=  -92896;
	5627: sound1 <=  -92224;
	5628: sound1 <=  -60608;
	5629: sound1 <=  -33356;
	5630: sound1 <=  -29602;
	5631: sound1 <=  -35736;
	5632: sound1 <=  -14984;
	5633: sound1 <=  57343;
	5634: sound1 <=  126770;
	5635: sound1 <=  202698;
	5636: sound1 <=  252716;
	5637: sound1 <=  271301;
	5638: sound1 <=  263855;
	5639: sound1 <=  241089;
	5640: sound1 <=  236328;
	5641: sound1 <=  280762;
	5642: sound1 <=  323334;
	5643: sound1 <=  324768;
	5644: sound1 <=  294586;
	5645: sound1 <=  275452;
	5646: sound1 <=  245667;
	5647: sound1 <=  247742;
	5648: sound1 <=  104187;
	5649: sound1 <=  -74951;
	5650: sound1 <=  -158661;
	5651: sound1 <=  -237732;
	5652: sound1 <=  -289886;
	5653: sound1 <=  -314362;
	5654: sound1 <=  -306458;
	5655: sound1 <=  -289642;
	5656: sound1 <=  -275513;
	5657: sound1 <=  -245300;
	5658: sound1 <=  -194061;
	5659: sound1 <=  -175110;
	5660: sound1 <=  -149719;
	5661: sound1 <=  -120911;
	5662: sound1 <=  -91034;
	5663: sound1 <=  -37750;
	5664: sound1 <=  13519;
	5665: sound1 <=  35583;
	5666: sound1 <=  48187;
	5667: sound1 <=  96649;
	5668: sound1 <=  131073;
	5669: sound1 <=  162933;
	5670: sound1 <=  220734;
	5671: sound1 <=  272552;
	5672: sound1 <=  177704;
	5673: sound1 <=  133972;
	5674: sound1 <=  160614;
	5675: sound1 <=  172913;
	5676: sound1 <=  199585;
	5677: sound1 <=  185699;
	5678: sound1 <=  174286;
	5679: sound1 <=  110962;
	5680: sound1 <=  46722;
	5681: sound1 <=  -71259;
	5682: sound1 <=  -230560;
	5683: sound1 <=  -251434;
	5684: sound1 <=  -274689;
	5685: sound1 <=  -275848;
	5686: sound1 <=  -283936;
	5687: sound1 <=  -259857;
	5688: sound1 <=  -262665;
	5689: sound1 <=  -272675;
	5690: sound1 <=  -281311;
	5691: sound1 <=  -288910;
	5692: sound1 <=  -267792;
	5693: sound1 <=  -231232;
	5694: sound1 <=  -185059;
	5695: sound1 <=  -126556;
	5696: sound1 <=  -66956;
	5697: sound1 <=  -12543;
	5698: sound1 <=  28534;
	5699: sound1 <=  89081;
	5700: sound1 <=  171936;
	5701: sound1 <=  210419;
	5702: sound1 <=  253235;
	5703: sound1 <=  314575;
	5704: sound1 <=  368530;
	5705: sound1 <=  372223;
	5706: sound1 <=  350555;
	5707: sound1 <=  318115;
	5708: sound1 <=  313904;
	5709: sound1 <=  320801;
	5710: sound1 <=  304108;
	5711: sound1 <=  305359;
	5712: sound1 <=  303955;
	5713: sound1 <=  327332;
	5714: sound1 <=  336792;
	5715: sound1 <=  337830;
	5716: sound1 <=  317139;
	5717: sound1 <=  307159;
	5718: sound1 <=  290161;
	5719: sound1 <=  263794;
	5720: sound1 <=  256500;
	5721: sound1 <=  232147;
	5722: sound1 <=  183167;
	5723: sound1 <=  145081;
	5724: sound1 <=  130646;
	5725: sound1 <=  106415;
	5726: sound1 <=  86700;
	5727: sound1 <=  76172;
	5728: sound1 <=  65460;
	5729: sound1 <=  41199;
	5730: sound1 <=  16602;
	5731: sound1 <=  30945;
	5732: sound1 <=  20996;
	5733: sound1 <=  -29327;
	5734: sound1 <=  -35339;
	5735: sound1 <=  -35858;
	5736: sound1 <=  -69244;
	5737: sound1 <=  -105591;
	5738: sound1 <=  -131683;
	5739: sound1 <=  -138428;
	5740: sound1 <=  -160767;
	5741: sound1 <=  -155365;
	5742: sound1 <=  -121948;
	5743: sound1 <=  -124023;
	5744: sound1 <=  -122620;
	5745: sound1 <=  -101654;
	5746: sound1 <=  -89600;
	5747: sound1 <=  -70160;
	5748: sound1 <=  -53650;
	5749: sound1 <=  -54474;
	5750: sound1 <=  -43427;
	5751: sound1 <=  -29999;
	5752: sound1 <=  -40466;
	5753: sound1 <=  -42969;
	5754: sound1 <=  -30090;
	5755: sound1 <=  -55969;
	5756: sound1 <=  -109589;
	5757: sound1 <=  -147552;
	5758: sound1 <=  -269592;
	5759: sound1 <=  -315918;
	5760: sound1 <=  -338409;
	5761: sound1 <=  -319489;
	5762: sound1 <=  -325867;
	5763: sound1 <=  -359894;
	5764: sound1 <=  -387268;
	5765: sound1 <=  -394257;
	5766: sound1 <=  -366913;
	5767: sound1 <=  -344604;
	5768: sound1 <=  -318939;
	5769: sound1 <=  -295288;
	5770: sound1 <=  -237518;
	5771: sound1 <=  -150146;
	5772: sound1 <=  -108063;
	5773: sound1 <=  -8423;
	5774: sound1 <=  79102;
	5775: sound1 <=  116058;
	5776: sound1 <=  163879;
	5777: sound1 <=  199219;
	5778: sound1 <=  212219;
	5779: sound1 <=  234772;
	5780: sound1 <=  241180;
	5781: sound1 <=  228210;
	5782: sound1 <=  203766;
	5783: sound1 <=  204437;
	5784: sound1 <=  240051;
	5785: sound1 <=  247772;
	5786: sound1 <=  243622;
	5787: sound1 <=  231720;
	5788: sound1 <=  215973;
	5789: sound1 <=  207184;
	5790: sound1 <=  204071;
	5791: sound1 <=  189301;
	5792: sound1 <=  184326;
	5793: sound1 <=  194824;
	5794: sound1 <=  192963;
	5795: sound1 <=  191742;
	5796: sound1 <=  180389;
	5797: sound1 <=  140747;
	5798: sound1 <=  112213;
	5799: sound1 <=  123688;
	5800: sound1 <=  132111;
	5801: sound1 <=  114655;
	5802: sound1 <=  119232;
	5803: sound1 <=  138000;
	5804: sound1 <=  144257;
	5805: sound1 <=  167755;
	5806: sound1 <=  174835;
	5807: sound1 <=  185272;
	5808: sound1 <=  195831;
	5809: sound1 <=  222992;
	5810: sound1 <=  286621;
	5811: sound1 <=  309265;
	5812: sound1 <=  296417;
	5813: sound1 <=  290588;
	5814: sound1 <=  303406;
	5815: sound1 <=  296692;
	5816: sound1 <=  277283;
	5817: sound1 <=  234192;
	5818: sound1 <=  163025;
	5819: sound1 <=  113190;
	5820: sound1 <=  90759;
	5821: sound1 <=  77759;
	5822: sound1 <=  23834;
	5823: sound1 <=  61;
	5824: sound1 <=  -14282;
	5825: sound1 <=  -14130;
	5826: sound1 <=  -28717;
	5827: sound1 <=  -23590;
	5828: sound1 <=  -14801;
	5829: sound1 <=  -1587;
	5830: sound1 <=  -9521;
	5831: sound1 <=  -43121;
	5832: sound1 <=  -60913;
	5833: sound1 <=  -89020;
	5834: sound1 <=  -97900;
	5835: sound1 <=  -110657;
	5836: sound1 <=  -135864;
	5837: sound1 <=  -224640;
	5838: sound1 <=  -360992;
	5839: sound1 <=  -347748;
	5840: sound1 <=  -336945;
	5841: sound1 <=  -351990;
	5842: sound1 <=  -372070;
	5843: sound1 <=  -363922;
	5844: sound1 <=  -370636;
	5845: sound1 <=  -371155;
	5846: sound1 <=  -351837;
	5847: sound1 <=  -359100;
	5848: sound1 <=  -352997;
	5849: sound1 <=  -354370;
	5850: sound1 <=  -371002;
	5851: sound1 <=  -334991;
	5852: sound1 <=  -279724;
	5853: sound1 <=  -212708;
	5854: sound1 <=  -179291;
	5855: sound1 <=  -202972;
	5856: sound1 <=  -153931;
	5857: sound1 <=  -156494;
	5858: sound1 <=  -106689;
	5859: sound1 <=  -35980;
	5860: sound1 <=  15167;
	5861: sound1 <=  84900;
	5862: sound1 <=  111786;
	5863: sound1 <=  132080;
	5864: sound1 <=  166321;
	5865: sound1 <=  166840;
	5866: sound1 <=  132080;
	5867: sound1 <=  87738;
	5868: sound1 <=  50507;
	5869: sound1 <=  26398;
	5870: sound1 <=  14862;
	5871: sound1 <=  -23102;
	5872: sound1 <=  -47211;
	5873: sound1 <=  -61493;
	5874: sound1 <=  -27374;
	5875: sound1 <=  17303;
	5876: sound1 <=  41840;
	5877: sound1 <=  56152;
	5878: sound1 <=  63141;
	5879: sound1 <=  26459;
	5880: sound1 <=  30426;
	5881: sound1 <=  64819;
	5882: sound1 <=  79773;
	5883: sound1 <=  73334;
	5884: sound1 <=  69244;
	5885: sound1 <=  97351;
	5886: sound1 <=  32990;
	5887: sound1 <=  47913;
	5888: sound1 <=  109680;
	5889: sound1 <=  63446;
	5890: sound1 <=  10803;
	5891: sound1 <=  53070;
	5892: sound1 <=  64972;
	5893: sound1 <=  124878;
	5894: sound1 <=  92346;
	5895: sound1 <=  111664;
	5896: sound1 <=  223236;
	5897: sound1 <=  210693;
	5898: sound1 <=  158234;
	5899: sound1 <=  194733;
	5900: sound1 <=  183533;
	5901: sound1 <=  210083;
	5902: sound1 <=  262054;
	5903: sound1 <=  193756;
	5904: sound1 <=  140594;
	5905: sound1 <=  115723;
	5906: sound1 <=  114105;
	5907: sound1 <=  150696;
	5908: sound1 <=  185211;
	5909: sound1 <=  234344;
	5910: sound1 <=  262939;
	5911: sound1 <=  285767;
	5912: sound1 <=  302185;
	5913: sound1 <=  289856;
	5914: sound1 <=  271210;
	5915: sound1 <=  236694;
	5916: sound1 <=  233185;
	5917: sound1 <=  97351;
	5918: sound1 <=  -4486;
	5919: sound1 <=  -39551;
	5920: sound1 <=  -101990;
	5921: sound1 <=  -129425;
	5922: sound1 <=  -140961;
	5923: sound1 <=  -138184;
	5924: sound1 <=  -102234;
	5925: sound1 <=  -62775;
	5926: sound1 <=  -54871;
	5927: sound1 <=  -43915;
	5928: sound1 <=  -9033;
	5929: sound1 <=  27863;
	5930: sound1 <=  87219;
	5931: sound1 <=  156036;
	5932: sound1 <=  210388;
	5933: sound1 <=  263306;
	5934: sound1 <=  319702;
	5935: sound1 <=  351013;
	5936: sound1 <=  362396;
	5937: sound1 <=  400208;
	5938: sound1 <=  431610;
	5939: sound1 <=  405914;
	5940: sound1 <=  390259;
	5941: sound1 <=  390015;
	5942: sound1 <=  370026;
	5943: sound1 <=  352020;
	5944: sound1 <=  306671;
	5945: sound1 <=  247650;
	5946: sound1 <=  235413;
	5947: sound1 <=  217651;
	5948: sound1 <=  165680;
	5949: sound1 <=  137238;
	5950: sound1 <=  98663;
	5951: sound1 <=  85785;
	5952: sound1 <=  56671;
	5953: sound1 <=  9338;
	5954: sound1 <=  -36865;
	5955: sound1 <=  -74341;
	5956: sound1 <=  -117523;
	5957: sound1 <=  -173309;
	5958: sound1 <=  -189423;
	5959: sound1 <=  -202423;
	5960: sound1 <=  -243439;
	5961: sound1 <=  -291626;
	5962: sound1 <=  -324738;
	5963: sound1 <=  -329132;
	5964: sound1 <=  -326141;
	5965: sound1 <=  -306519;
	5966: sound1 <=  -278229;
	5967: sound1 <=  -208466;
	5968: sound1 <=  -157745;
	5969: sound1 <=  -113251;
	5970: sound1 <=  -80475;
	5971: sound1 <=  -80261;
	5972: sound1 <=  -85144;
	5973: sound1 <=  -100464;
	5974: sound1 <=  -94543;
	5975: sound1 <=  -56702;
	5976: sound1 <=  -44495;
	5977: sound1 <=  -29144;
	5978: sound1 <=  -54749;
	5979: sound1 <=  -83374;
	5980: sound1 <=  -88104;
	5981: sound1 <=  -96100;
	5982: sound1 <=  -100647;
	5983: sound1 <=  -118652;
	5984: sound1 <=  -143066;
	5985: sound1 <=  -184296;
	5986: sound1 <=  -182861;
	5987: sound1 <=  -165192;
	5988: sound1 <=  -149078;
	5989: sound1 <=  -152161;
	5990: sound1 <=  -112549;
	5991: sound1 <=  -65765;
	5992: sound1 <=  -15656;
	5993: sound1 <=  51086;
	5994: sound1 <=  126190;
	5995: sound1 <=  172729;
	5996: sound1 <=  173615;
	5997: sound1 <=  153168;
	5998: sound1 <=  161255;
	5999: sound1 <=  179565;
	6000: sound1 <=  198334;
	6001: sound1 <=  203430;
	6002: sound1 <=  180786;
	6003: sound1 <=  157074;
	6004: sound1 <=  141998;
	6005: sound1 <=  123535;
	6006: sound1 <=  101196;
	6007: sound1 <=  73425;
	6008: sound1 <=  76111;
	6009: sound1 <=  56824;
	6010: sound1 <=  15839;
	6011: sound1 <=  15717;
	6012: sound1 <=  34393;
	6013: sound1 <=  23743;
	6014: sound1 <=  -20752;
	6015: sound1 <=  -23346;
	6016: sound1 <=  -11749;
	6017: sound1 <=  -20142;
	6018: sound1 <=  -3418;
	6019: sound1 <=  -61707;
	6020: sound1 <=  -167236;
	6021: sound1 <=  -185089;
	6022: sound1 <=  -228851;
	6023: sound1 <=  -275513;
	6024: sound1 <=  -303040;
	6025: sound1 <=  -275848;
	6026: sound1 <=  -263885;
	6027: sound1 <=  -228577;
	6028: sound1 <=  -172791;
	6029: sound1 <=  -134827;
	6030: sound1 <=  -91980;
	6031: sound1 <=  -54962;
	6032: sound1 <=  -32745;
	6033: sound1 <=  13702;
	6034: sound1 <=  111877;
	6035: sound1 <=  188385;
	6036: sound1 <=  238800;
	6037: sound1 <=  299713;
	6038: sound1 <=  337067;
	6039: sound1 <=  359894;
	6040: sound1 <=  359131;
	6041: sound1 <=  346313;
	6042: sound1 <=  363983;
	6043: sound1 <=  352814;
	6044: sound1 <=  328033;
	6045: sound1 <=  311829;
	6046: sound1 <=  299011;
	6047: sound1 <=  300598;
	6048: sound1 <=  300720;
	6049: sound1 <=  278992;
	6050: sound1 <=  257477;
	6051: sound1 <=  246582;
	6052: sound1 <=  238953;
	6053: sound1 <=  224487;
	6054: sound1 <=  196106;
	6055: sound1 <=  164886;
	6056: sound1 <=  150482;
	6057: sound1 <=  107697;
	6058: sound1 <=  92621;
	6059: sound1 <=  87158;
	6060: sound1 <=  72357;
	6061: sound1 <=  93018;
	6062: sound1 <=  140350;
	6063: sound1 <=  145569;
	6064: sound1 <=  125275;
	6065: sound1 <=  74493;
	6066: sound1 <=  62286;
	6067: sound1 <=  48798;
	6068: sound1 <=  41931;
	6069: sound1 <=  15350;
	6070: sound1 <=  -22552;
	6071: sound1 <=  14343;
	6072: sound1 <=  22003;
	6073: sound1 <=  25146;
	6074: sound1 <=  27649;
	6075: sound1 <=  3052;
	6076: sound1 <=  -16266;
	6077: sound1 <=  -44403;
	6078: sound1 <=  -122467;
	6079: sound1 <=  -174835;
	6080: sound1 <=  -200409;
	6081: sound1 <=  -234863;
	6082: sound1 <=  -234497;
	6083: sound1 <=  -236786;
	6084: sound1 <=  -259796;
	6085: sound1 <=  -279846;
	6086: sound1 <=  -289063;
	6087: sound1 <=  -282104;
	6088: sound1 <=  -275146;
	6089: sound1 <=  -298096;
	6090: sound1 <=  -335785;
	6091: sound1 <=  -353607;
	6092: sound1 <=  -358368;
	6093: sound1 <=  -332397;
	6094: sound1 <=  -290863;
	6095: sound1 <=  -262665;
	6096: sound1 <=  -249512;
	6097: sound1 <=  -224304;
	6098: sound1 <=  -178406;
	6099: sound1 <=  -127167;
	6100: sound1 <=  -99457;
	6101: sound1 <=  -84595;
	6102: sound1 <=  -73090;
	6103: sound1 <=  -56549;
	6104: sound1 <=  -21576;
	6105: sound1 <=  18005;
	6106: sound1 <=  49622;
	6107: sound1 <=  67627;
	6108: sound1 <=  99976;
	6109: sound1 <=  147034;
	6110: sound1 <=  158112;
	6111: sound1 <=  169434;
	6112: sound1 <=  166107;
	6113: sound1 <=  117279;
	6114: sound1 <=  102325;
	6115: sound1 <=  125946;
	6116: sound1 <=  154144;
	6117: sound1 <=  163086;
	6118: sound1 <=  168732;
	6119: sound1 <=  205139;
	6120: sound1 <=  222076;
	6121: sound1 <=  231689;
	6122: sound1 <=  212158;
	6123: sound1 <=  207672;
	6124: sound1 <=  204712;
	6125: sound1 <=  201477;
	6126: sound1 <=  190338;
	6127: sound1 <=  148102;
	6128: sound1 <=  138031;
	6129: sound1 <=  142456;
	6130: sound1 <=  111969;
	6131: sound1 <=  92560;
	6132: sound1 <=  89691;
	6133: sound1 <=  78644;
	6134: sound1 <=  42725;
	6135: sound1 <=  -109222;
	6136: sound1 <=  -98907;
	6137: sound1 <=  -48584;
	6138: sound1 <=  -74402;
	6139: sound1 <=  -113525;
	6140: sound1 <=  -98694;
	6141: sound1 <=  -98633;
	6142: sound1 <=  -59631;
	6143: sound1 <=  -22797;
	6144: sound1 <=  -31;
	6145: sound1 <=  26825;
	6146: sound1 <=  56244;
	6147: sound1 <=  101532;
	6148: sound1 <=  154358;
	6149: sound1 <=  227936;
	6150: sound1 <=  215729;
	6151: sound1 <=  203583;
	6152: sound1 <=  236664;
	6153: sound1 <=  221008;
	6154: sound1 <=  211060;
	6155: sound1 <=  199707;
	6156: sound1 <=  169800;
	6157: sound1 <=  156128;
	6158: sound1 <=  180908;
	6159: sound1 <=  186371;
	6160: sound1 <=  204895;
	6161: sound1 <=  199585;
	6162: sound1 <=  193451;
	6163: sound1 <=  77911;
	6164: sound1 <=  47974;
	6165: sound1 <=  77423;
	6166: sound1 <=  77271;
	6167: sound1 <=  78217;
	6168: sound1 <=  71442;
	6169: sound1 <=  88440;
	6170: sound1 <=  73242;
	6171: sound1 <=  50079;
	6172: sound1 <=  45044;
	6173: sound1 <=  29968;
	6174: sound1 <=  -57648;
	6175: sound1 <=  -186340;
	6176: sound1 <=  -215729;
	6177: sound1 <=  -226807;
	6178: sound1 <=  -206604;
	6179: sound1 <=  -187592;
	6180: sound1 <=  -203461;
	6181: sound1 <=  -220032;
	6182: sound1 <=  -189240;
	6183: sound1 <=  -154114;
	6184: sound1 <=  -100952;
	6185: sound1 <=  -53253;
	6186: sound1 <=  -21088;
	6187: sound1 <=  27893;
	6188: sound1 <=  56824;
	6189: sound1 <=  56824;
	6190: sound1 <=  70496;
	6191: sound1 <=  120514;
	6192: sound1 <=  174103;
	6193: sound1 <=  201691;
	6194: sound1 <=  197113;
	6195: sound1 <=  192108;
	6196: sound1 <=  196564;
	6197: sound1 <=  199860;
	6198: sound1 <=  218353;
	6199: sound1 <=  244354;
	6200: sound1 <=  259399;
	6201: sound1 <=  272583;
	6202: sound1 <=  287720;
	6203: sound1 <=  278961;
	6204: sound1 <=  279083;
	6205: sound1 <=  287445;
	6206: sound1 <=  275330;
	6207: sound1 <=  234406;
	6208: sound1 <=  200989;
	6209: sound1 <=  152954;
	6210: sound1 <=  107513;
	6211: sound1 <=  74219;
	6212: sound1 <=  64209;
	6213: sound1 <=  73456;
	6214: sound1 <=  72968;
	6215: sound1 <=  99091;
	6216: sound1 <=  -27435;
	6217: sound1 <=  -101685;
	6218: sound1 <=  -97565;
	6219: sound1 <=  -107483;
	6220: sound1 <=  -88867;
	6221: sound1 <=  -73761;
	6222: sound1 <=  -52032;
	6223: sound1 <=  -81238;
	6224: sound1 <=  -125793;
	6225: sound1 <=  -127380;
	6226: sound1 <=  -104156;
	6227: sound1 <=  -87860;
	6228: sound1 <=  -62408;
	6229: sound1 <=  -72937;
	6230: sound1 <=  -73853;
	6231: sound1 <=  -36102;
	6232: sound1 <=  10620;
	6233: sound1 <=  50720;
	6234: sound1 <=  91736;
	6235: sound1 <=  106140;
	6236: sound1 <=  98724;
	6237: sound1 <=  111725;
	6238: sound1 <=  91522;
	6239: sound1 <=  122406;
	6240: sound1 <=  27496;
	6241: sound1 <=  -103729;
	6242: sound1 <=  -107971;
	6243: sound1 <=  -162842;
	6244: sound1 <=  -217712;
	6245: sound1 <=  -278381;
	6246: sound1 <=  -285583;
	6247: sound1 <=  -290680;
	6248: sound1 <=  -304321;
	6249: sound1 <=  -316772;
	6250: sound1 <=  -323212;
	6251: sound1 <=  -319397;
	6252: sound1 <=  -256317;
	6253: sound1 <=  -176239;
	6254: sound1 <=  -125732;
	6255: sound1 <=  -78339;
	6256: sound1 <=  -60852;
	6257: sound1 <=  -22736;
	6258: sound1 <=  10193;
	6259: sound1 <=  46387;
	6260: sound1 <=  57312;
	6261: sound1 <=  81635;
	6262: sound1 <=  112457;
	6263: sound1 <=  164398;
	6264: sound1 <=  226715;
	6265: sound1 <=  271606;
	6266: sound1 <=  281769;
	6267: sound1 <=  292969;
	6268: sound1 <=  309937;
	6269: sound1 <=  290161;
	6270: sound1 <=  269989;
	6271: sound1 <=  280457;
	6272: sound1 <=  274750;
	6273: sound1 <=  268707;
	6274: sound1 <=  287872;
	6275: sound1 <=  284149;
	6276: sound1 <=  284790;
	6277: sound1 <=  263245;
	6278: sound1 <=  230225;
	6279: sound1 <=  225952;
	6280: sound1 <=  218842;
	6281: sound1 <=  209167;
	6282: sound1 <=  205780;
	6283: sound1 <=  184784;
	6284: sound1 <=  152863;
	6285: sound1 <=  142365;
	6286: sound1 <=  97717;
	6287: sound1 <=  65216;
	6288: sound1 <=  35278;
	6289: sound1 <=  8545;
	6290: sound1 <=  18707;
	6291: sound1 <=  49316;
	6292: sound1 <=  81177;
	6293: sound1 <=  105438;
	6294: sound1 <=  108429;
	6295: sound1 <=  100311;
	6296: sound1 <=  80566;
	6297: sound1 <=  86395;
	6298: sound1 <=  80322;
	6299: sound1 <=  57312;
	6300: sound1 <=  36713;
	6301: sound1 <=  26855;
	6302: sound1 <=  16663;
	6303: sound1 <=  7538;
	6304: sound1 <=  -8942;
	6305: sound1 <=  -41290;
	6306: sound1 <=  -70251;
	6307: sound1 <=  -110138;
	6308: sound1 <=  -152252;
	6309: sound1 <=  -175293;
	6310: sound1 <=  -184082;
	6311: sound1 <=  -198730;
	6312: sound1 <=  -236725;
	6313: sound1 <=  -270111;
	6314: sound1 <=  -288666;
	6315: sound1 <=  -353424;
	6316: sound1 <=  -383423;
	6317: sound1 <=  -367584;
	6318: sound1 <=  -361786;
	6319: sound1 <=  -394226;
	6320: sound1 <=  -408844;
	6321: sound1 <=  -410309;
	6322: sound1 <=  -398651;
	6323: sound1 <=  -376495;
	6324: sound1 <=  -326843;
	6325: sound1 <=  -256348;
	6326: sound1 <=  -203522;
	6327: sound1 <=  -149384;
	6328: sound1 <=  -55389;
	6329: sound1 <=  11536;
	6330: sound1 <=  -52795;
	6331: sound1 <=  -24384;
	6332: sound1 <=  57526;
	6333: sound1 <=  134338;
	6334: sound1 <=  204773;
	6335: sound1 <=  189331;
	6336: sound1 <=  193054;
	6337: sound1 <=  191681;
	6338: sound1 <=  174713;
	6339: sound1 <=  134338;
	6340: sound1 <=  130646;
	6341: sound1 <=  110260;
	6342: sound1 <=  120758;
	6343: sound1 <=  72083;
	6344: sound1 <=  89203;
	6345: sound1 <=  138000;
	6346: sound1 <=  85510;
	6347: sound1 <=  21149;
	6348: sound1 <=  43945;
	6349: sound1 <=  31891;
	6350: sound1 <=  -65369;
	6351: sound1 <=  -62988;
	6352: sound1 <=  -47272;
	6353: sound1 <=  -114014;
	6354: sound1 <=  -78644;
	6355: sound1 <=  -101776;
	6356: sound1 <=  -98083;
	6357: sound1 <=  -40558;
	6358: sound1 <=  -28900;
	6359: sound1 <=  -22705;
	6360: sound1 <=  -183;
	6361: sound1 <=  -17151;
	6362: sound1 <=  -27405;
	6363: sound1 <=  16357;
	6364: sound1 <=  67688;
	6365: sound1 <=  33020;
	6366: sound1 <=  -5219;
	6367: sound1 <=  54993;
	6368: sound1 <=  74585;
	6369: sound1 <=  102936;
	6370: sound1 <=  60364;
	6371: sound1 <=  143738;
	6372: sound1 <=  126892;
	6373: sound1 <=  85541;
	6374: sound1 <=  151428;
	6375: sound1 <=  81116;
	6376: sound1 <=  81055;
	6377: sound1 <=  131836;
	6378: sound1 <=  141876;
	6379: sound1 <=  155792;
	6380: sound1 <=  116821;
	6381: sound1 <=  27100;
	6382: sound1 <=  50507;
	6383: sound1 <=  61401;
	6384: sound1 <=  66223;
	6385: sound1 <=  81146;
	6386: sound1 <=  101837;
	6387: sound1 <=  89966;
	6388: sound1 <=  -3418;
	6389: sound1 <=  -16754;
	6390: sound1 <=  24475;
	6391: sound1 <=  55786;
	6392: sound1 <=  58197;
	6393: sound1 <=  92102;
	6394: sound1 <=  121765;
	6395: sound1 <=  127808;
	6396: sound1 <=  119415;
	6397: sound1 <=  95032;
	6398: sound1 <=  101013;
	6399: sound1 <=  145874;
	6400: sound1 <=  148041;
	6401: sound1 <=  173157;
	6402: sound1 <=  182434;
	6403: sound1 <=  163940;
	6404: sound1 <=  161285;
	6405: sound1 <=  169403;
	6406: sound1 <=  156128;
	6407: sound1 <=  143677;
	6408: sound1 <=  128632;
	6409: sound1 <=  123413;
	6410: sound1 <=  134094;
	6411: sound1 <=  134155;
	6412: sound1 <=  133301;
	6413: sound1 <=  144226;
	6414: sound1 <=  131805;
	6415: sound1 <=  102509;
	6416: sound1 <=  77942;
	6417: sound1 <=  87402;
	6418: sound1 <=  61066;
	6419: sound1 <=  30243;
	6420: sound1 <=  22522;
	6421: sound1 <=  24506;
	6422: sound1 <=  29053;
	6423: sound1 <=  34607;
	6424: sound1 <=  53833;
	6425: sound1 <=  73761;
	6426: sound1 <=  74188;
	6427: sound1 <=  -33722;
	6428: sound1 <=  -110626;
	6429: sound1 <=  -128723;
	6430: sound1 <=  -179688;
	6431: sound1 <=  -210052;
	6432: sound1 <=  -206116;
	6433: sound1 <=  -193939;
	6434: sound1 <=  -197845;
	6435: sound1 <=  -226868;
	6436: sound1 <=  -249359;
	6437: sound1 <=  -232513;
	6438: sound1 <=  -182190;
	6439: sound1 <=  -126587;
	6440: sound1 <=  -89417;
	6441: sound1 <=  -45868;
	6442: sound1 <=  92;
	6443: sound1 <=  30273;
	6444: sound1 <=  51575;
	6445: sound1 <=  67108;
	6446: sound1 <=  83282;
	6447: sound1 <=  112793;
	6448: sound1 <=  142822;
	6449: sound1 <=  182068;
	6450: sound1 <=  215912;
	6451: sound1 <=  234344;
	6452: sound1 <=  250153;
	6453: sound1 <=  278015;
	6454: sound1 <=  312744;
	6455: sound1 <=  310333;
	6456: sound1 <=  308258;
	6457: sound1 <=  308929;
	6458: sound1 <=  339508;
	6459: sound1 <=  382324;
	6460: sound1 <=  387054;
	6461: sound1 <=  392487;
	6462: sound1 <=  379669;
	6463: sound1 <=  349518;
	6464: sound1 <=  325684;
	6465: sound1 <=  301819;
	6466: sound1 <=  259155;
	6467: sound1 <=  237976;
	6468: sound1 <=  236908;
	6469: sound1 <=  232269;
	6470: sound1 <=  237366;
	6471: sound1 <=  207428;
	6472: sound1 <=  190765;
	6473: sound1 <=  170563;
	6474: sound1 <=  164215;
	6475: sound1 <=  133362;
	6476: sound1 <=  72510;
	6477: sound1 <=  7324;
	6478: sound1 <=  -51788;
	6479: sound1 <=  -84656;
	6480: sound1 <=  -115417;
	6481: sound1 <=  -155579;
	6482: sound1 <=  -206543;
	6483: sound1 <=  -226013;
	6484: sound1 <=  -258820;
	6485: sound1 <=  -252350;
	6486: sound1 <=  -254120;
	6487: sound1 <=  -258759;
	6488: sound1 <=  -226044;
	6489: sound1 <=  -204742;
	6490: sound1 <=  -227203;
	6491: sound1 <=  -254150;
	6492: sound1 <=  -253082;
	6493: sound1 <=  -235809;
	6494: sound1 <=  -211670;
	6495: sound1 <=  -218994;
	6496: sound1 <=  -236816;
	6497: sound1 <=  -242889;
	6498: sound1 <=  -242004;
	6499: sound1 <=  -238556;
	6500: sound1 <=  -218903;
	6501: sound1 <=  -214417;
	6502: sound1 <=  -213623;
	6503: sound1 <=  -202057;
	6504: sound1 <=  -202667;
	6505: sound1 <=  -196960;
	6506: sound1 <=  -204742;
	6507: sound1 <=  -221100;
	6508: sound1 <=  -231720;
	6509: sound1 <=  -216858;
	6510: sound1 <=  -209351;
	6511: sound1 <=  -196472;
	6512: sound1 <=  -179443;
	6513: sound1 <=  -155029;
	6514: sound1 <=  -121948;
	6515: sound1 <=  -95551;
	6516: sound1 <=  -62378;
	6517: sound1 <=  -23010;
	6518: sound1 <=  -366;
	6519: sound1 <=  3540;
	6520: sound1 <=  8545;
	6521: sound1 <=  56763;
	6522: sound1 <=  101074;
	6523: sound1 <=  115143;
	6524: sound1 <=  137543;
	6525: sound1 <=  141449;
	6526: sound1 <=  129333;
	6527: sound1 <=  135468;
	6528: sound1 <=  140930;
	6529: sound1 <=  155487;
	6530: sound1 <=  181732;
	6531: sound1 <=  183075;
	6532: sound1 <=  31067;
	6533: sound1 <=  -29663;
	6534: sound1 <=  -34454;
	6535: sound1 <=  -75073;
	6536: sound1 <=  -98785;
	6537: sound1 <=  -103088;
	6538: sound1 <=  -89691;
	6539: sound1 <=  -124542;
	6540: sound1 <=  -137573;
	6541: sound1 <=  -86090;
	6542: sound1 <=  -23529;
	6543: sound1 <=  37506;
	6544: sound1 <=  89264;
	6545: sound1 <=  154144;
	6546: sound1 <=  203888;
	6547: sound1 <=  229279;
	6548: sound1 <=  247772;
	6549: sound1 <=  291016;
	6550: sound1 <=  313599;
	6551: sound1 <=  326172;
	6552: sound1 <=  346497;
	6553: sound1 <=  369629;
	6554: sound1 <=  383972;
	6555: sound1 <=  393707;
	6556: sound1 <=  418854;
	6557: sound1 <=  441711;
	6558: sound1 <=  448883;
	6559: sound1 <=  440460;
	6560: sound1 <=  419312;
	6561: sound1 <=  403259;
	6562: sound1 <=  405670;
	6563: sound1 <=  407562;
	6564: sound1 <=  419434;
	6565: sound1 <=  409546;
	6566: sound1 <=  399536;
	6567: sound1 <=  365631;
	6568: sound1 <=  313660;
	6569: sound1 <=  300629;
	6570: sound1 <=  266266;
	6571: sound1 <=  214569;
	6572: sound1 <=  164215;
	6573: sound1 <=  112610;
	6574: sound1 <=  75989;
	6575: sound1 <=  42633;
	6576: sound1 <=  -7355;
	6577: sound1 <=  -69427;
	6578: sound1 <=  -115082;
	6579: sound1 <=  -165680;
	6580: sound1 <=  -190613;
	6581: sound1 <=  -178741;
	6582: sound1 <=  -185120;
	6583: sound1 <=  -159180;
	6584: sound1 <=  -121674;
	6585: sound1 <=  -118896;
	6586: sound1 <=  -105194;
	6587: sound1 <=  -99579;
	6588: sound1 <=  -92438;
	6589: sound1 <=  -90485;
	6590: sound1 <=  -109985;
	6591: sound1 <=  -133911;
	6592: sound1 <=  -124084;
	6593: sound1 <=  -129059;
	6594: sound1 <=  -157837;
	6595: sound1 <=  -153656;
	6596: sound1 <=  -152435;
	6597: sound1 <=  -142517;
	6598: sound1 <=  -158813;
	6599: sound1 <=  -172882;
	6600: sound1 <=  -186859;
	6601: sound1 <=  -177216;
	6602: sound1 <=  -225372;
	6603: sound1 <=  -306488;
	6604: sound1 <=  -300018;
	6605: sound1 <=  -288391;
	6606: sound1 <=  -286743;
	6607: sound1 <=  -294128;
	6608: sound1 <=  -292694;
	6609: sound1 <=  -300598;
	6610: sound1 <=  -286774;
	6611: sound1 <=  -263245;
	6612: sound1 <=  -190918;
	6613: sound1 <=  -114716;
	6614: sound1 <=  -81635;
	6615: sound1 <=  -55908;
	6616: sound1 <=  -49469;
	6617: sound1 <=  -143829;
	6618: sound1 <=  -109619;
	6619: sound1 <=  -48553;
	6620: sound1 <=  -10132;
	6621: sound1 <=  28046;
	6622: sound1 <=  32745;
	6623: sound1 <=  38635;
	6624: sound1 <=  62714;
	6625: sound1 <=  78827;
	6626: sound1 <=  124847;
	6627: sound1 <=  167908;
	6628: sound1 <=  194763;
	6629: sound1 <=  209900;
	6630: sound1 <=  235992;
	6631: sound1 <=  299561;
	6632: sound1 <=  309265;
	6633: sound1 <=  328094;
	6634: sound1 <=  279633;
	6635: sound1 <=  200836;
	6636: sound1 <=  187683;
	6637: sound1 <=  115753;
	6638: sound1 <=  98816;
	6639: sound1 <=  128784;
	6640: sound1 <=  173737;
	6641: sound1 <=  218933;
	6642: sound1 <=  220764;
	6643: sound1 <=  201965;
	6644: sound1 <=  184998;
	6645: sound1 <=  181824;
	6646: sound1 <=  169403;
	6647: sound1 <=  117920;
	6648: sound1 <=  -58533;
	6649: sound1 <=  -139465;
	6650: sound1 <=  -143127;
	6651: sound1 <=  -102539;
	6652: sound1 <=  -44739;
	6653: sound1 <=  3662;
	6654: sound1 <=  62500;
	6655: sound1 <=  82367;
	6656: sound1 <=  74646;
	6657: sound1 <=  82153;
	6658: sound1 <=  87555;
	6659: sound1 <=  91217;
	6660: sound1 <=  128143;
	6661: sound1 <=  163574;
	6662: sound1 <=  156219;
	6663: sound1 <=  146820;
	6664: sound1 <=  122681;
	6665: sound1 <=  108826;
	6666: sound1 <=  72754;
	6667: sound1 <=  -42358;
	6668: sound1 <=  -55939;
	6669: sound1 <=  -89050;
	6670: sound1 <=  -105896;
	6671: sound1 <=  -96832;
	6672: sound1 <=  -80353;
	6673: sound1 <=  -33905;
	6674: sound1 <=  18127;
	6675: sound1 <=  80292;
	6676: sound1 <=  146637;
	6677: sound1 <=  160950;
	6678: sound1 <=  185425;
	6679: sound1 <=  111633;
	6680: sound1 <=  -28412;
	6681: sound1 <=  -50476;
	6682: sound1 <=  -83862;
	6683: sound1 <=  -105194;
	6684: sound1 <=  -147461;
	6685: sound1 <=  -183746;
	6686: sound1 <=  -145294;
	6687: sound1 <=  -109680;
	6688: sound1 <=  -88226;
	6689: sound1 <=  -45959;
	6690: sound1 <=  -6500;
	6691: sound1 <=  29510;
	6692: sound1 <=  86060;
	6693: sound1 <=  144257;
	6694: sound1 <=  161865;
	6695: sound1 <=  188751;
	6696: sound1 <=  228088;
	6697: sound1 <=  258453;
	6698: sound1 <=  286926;
	6699: sound1 <=  331940;
	6700: sound1 <=  350342;
	6701: sound1 <=  350952;
	6702: sound1 <=  346252;
	6703: sound1 <=  334015;
	6704: sound1 <=  306396;
	6705: sound1 <=  270691;
	6706: sound1 <=  245972;
	6707: sound1 <=  254395;
	6708: sound1 <=  251556;
	6709: sound1 <=  227448;
	6710: sound1 <=  78918;
	6711: sound1 <=  -1465;
	6712: sound1 <=  -73212;
	6713: sound1 <=  -149292;
	6714: sound1 <=  -204956;
	6715: sound1 <=  -249664;
	6716: sound1 <=  -272278;
	6717: sound1 <=  -286865;
	6718: sound1 <=  -303711;
	6719: sound1 <=  -290833;
	6720: sound1 <=  -264648;
	6721: sound1 <=  -244232;
	6722: sound1 <=  -240967;
	6723: sound1 <=  -214874;
	6724: sound1 <=  -151367;
	6725: sound1 <=  -79529;
	6726: sound1 <=  -23102;
	6727: sound1 <=  12573;
	6728: sound1 <=  63324;
	6729: sound1 <=  96436;
	6730: sound1 <=  110229;
	6731: sound1 <=  155701;
	6732: sound1 <=  125702;
	6733: sound1 <=  130371;
	6734: sound1 <=  177063;
	6735: sound1 <=  207825;
	6736: sound1 <=  207275;
	6737: sound1 <=  199493;
	6738: sound1 <=  167511;
	6739: sound1 <=  149384;
	6740: sound1 <=  78339;
	6741: sound1 <=  -29755;
	6742: sound1 <=  -34302;
	6743: sound1 <=  -30212;
	6744: sound1 <=  4181;
	6745: sound1 <=  -45959;
	6746: sound1 <=  -127655;
	6747: sound1 <=  -112885;
	6748: sound1 <=  -96619;
	6749: sound1 <=  -149323;
	6750: sound1 <=  -183472;
	6751: sound1 <=  -110687;
	6752: sound1 <=  -149841;
	6753: sound1 <=  -223389;
	6754: sound1 <=  -165222;
	6755: sound1 <=  -87402;
	6756: sound1 <=  -125824;
	6757: sound1 <=  -86365;
	6758: sound1 <=  -55511;
	6759: sound1 <=  -31830;
	6760: sound1 <=  1099;
	6761: sound1 <=  5005;
	6762: sound1 <=  7538;
	6763: sound1 <=  -2899;
	6764: sound1 <=  -20508;
	6765: sound1 <=  -24902;
	6766: sound1 <=  29236;
	6767: sound1 <=  66895;
	6768: sound1 <=  75439;
	6769: sound1 <=  89844;
	6770: sound1 <=  82977;
	6771: sound1 <=  52734;
	6772: sound1 <=  33081;
	6773: sound1 <=  13306;
	6774: sound1 <=  36407;
	6775: sound1 <=  25482;
	6776: sound1 <=  -2472;
	6777: sound1 <=  -24536;
	6778: sound1 <=  12360;
	6779: sound1 <=  3021;
	6780: sound1 <=  -2075;
	6781: sound1 <=  -36194;
	6782: sound1 <=  -17761;
	6783: sound1 <=  -15869;
	6784: sound1 <=  12299;
	6785: sound1 <=  26947;
	6786: sound1 <=  -22247;
	6787: sound1 <=  18677;
	6788: sound1 <=  26581;
	6789: sound1 <=  -31219;
	6790: sound1 <=  3082;
	6791: sound1 <=  32349;
	6792: sound1 <=  46814;
	6793: sound1 <=  -50079;
	6794: sound1 <=  -95673;
	6795: sound1 <=  -106720;
	6796: sound1 <=  -81787;
	6797: sound1 <=  -14069;
	6798: sound1 <=  18921;
	6799: sound1 <=  49377;
	6800: sound1 <=  92468;
	6801: sound1 <=  139191;
	6802: sound1 <=  171082;
	6803: sound1 <=  184448;
	6804: sound1 <=  201416;
	6805: sound1 <=  97473;
	6806: sound1 <=  73120;
	6807: sound1 <=  109131;
	6808: sound1 <=  121674;
	6809: sound1 <=  120026;
	6810: sound1 <=  123840;
	6811: sound1 <=  133606;
	6812: sound1 <=  161926;
	6813: sound1 <=  186493;
	6814: sound1 <=  199097;
	6815: sound1 <=  203003;
	6816: sound1 <=  205078;
	6817: sound1 <=  205566;
	6818: sound1 <=  215027;
	6819: sound1 <=  226471;
	6820: sound1 <=  233734;
	6821: sound1 <=  200623;
	6822: sound1 <=  70770;
	6823: sound1 <=  21332;
	6824: sound1 <=  9216;
	6825: sound1 <=  -4211;
	6826: sound1 <=  -13489;
	6827: sound1 <=  -17120;
	6828: sound1 <=  -16876;
	6829: sound1 <=  -20782;
	6830: sound1 <=  -39368;
	6831: sound1 <=  -59967;
	6832: sound1 <=  -29358;
	6833: sound1 <=  732;
	6834: sound1 <=  8057;
	6835: sound1 <=  19073;
	6836: sound1 <=  13184;
	6837: sound1 <=  39825;
	6838: sound1 <=  84076;
	6839: sound1 <=  102264;
	6840: sound1 <=  154236;
	6841: sound1 <=  165039;
	6842: sound1 <=  168945;
	6843: sound1 <=  184357;
	6844: sound1 <=  217041;
	6845: sound1 <=  249298;
	6846: sound1 <=  281982;
	6847: sound1 <=  282623;
	6848: sound1 <=  268127;
	6849: sound1 <=  243744;
	6850: sound1 <=  219147;
	6851: sound1 <=  226715;
	6852: sound1 <=  232635;
	6853: sound1 <=  222321;
	6854: sound1 <=  218842;
	6855: sound1 <=  201233;
	6856: sound1 <=  203369;
	6857: sound1 <=  210754;
	6858: sound1 <=  162903;
	6859: sound1 <=  152557;
	6860: sound1 <=  169281;
	6861: sound1 <=  162476;
	6862: sound1 <=  126099;
	6863: sound1 <=  126770;
	6864: sound1 <=  105438;
	6865: sound1 <=  75775;
	6866: sound1 <=  54810;
	6867: sound1 <=  19623;
	6868: sound1 <=  -27588;
	6869: sound1 <=  -75500;
	6870: sound1 <=  -91400;
	6871: sound1 <=  -88715;
	6872: sound1 <=  -88898;
	6873: sound1 <=  -107635;
	6874: sound1 <=  -118317;
	6875: sound1 <=  -145081;
	6876: sound1 <=  -173981;
	6877: sound1 <=  -195282;
	6878: sound1 <=  -219727;
	6879: sound1 <=  -233551;
	6880: sound1 <=  -242676;
	6881: sound1 <=  -236206;
	6882: sound1 <=  -230560;
	6883: sound1 <=  -224457;
	6884: sound1 <=  -213074;
	6885: sound1 <=  -206970;
	6886: sound1 <=  -218079;
	6887: sound1 <=  -234589;
	6888: sound1 <=  -247650;
	6889: sound1 <=  -271637;
	6890: sound1 <=  -293304;
	6891: sound1 <=  -302521;
	6892: sound1 <=  -274139;
	6893: sound1 <=  -258606;
	6894: sound1 <=  -262238;
	6895: sound1 <=  -264130;
	6896: sound1 <=  -263000;
	6897: sound1 <=  -256744;
	6898: sound1 <=  -253540;
	6899: sound1 <=  -245728;
	6900: sound1 <=  -241455;
	6901: sound1 <=  -240204;
	6902: sound1 <=  -211639;
	6903: sound1 <=  -150177;
	6904: sound1 <=  -111603;
	6905: sound1 <=  -44800;
	6906: sound1 <=  -2472;
	6907: sound1 <=  60730;
	6908: sound1 <=  109161;
	6909: sound1 <=  128784;
	6910: sound1 <=  163147;
	6911: sound1 <=  192657;
	6912: sound1 <=  206390;
	6913: sound1 <=  233917;
	6914: sound1 <=  239075;
	6915: sound1 <=  214722;
	6916: sound1 <=  222473;
	6917: sound1 <=  250305;
	6918: sound1 <=  293335;
	6919: sound1 <=  285156;
	6920: sound1 <=  245117;
	6921: sound1 <=  203522;
	6922: sound1 <=  204376;
	6923: sound1 <=  220764;
	6924: sound1 <=  226624;
	6925: sound1 <=  189728;
	6926: sound1 <=  182251;
	6927: sound1 <=  206360;
	6928: sound1 <=  209991;
	6929: sound1 <=  211823;
	6930: sound1 <=  186523;
	6931: sound1 <=  167511;
	6932: sound1 <=  168427;
	6933: sound1 <=  177032;
	6934: sound1 <=  194611;
	6935: sound1 <=  197906;
	6936: sound1 <=  193207;
	6937: sound1 <=  199585;
	6938: sound1 <=  181488;
	6939: sound1 <=  159882;
	6940: sound1 <=  169312;
	6941: sound1 <=  173584;
	6942: sound1 <=  156616;
	6943: sound1 <=  141785;
	6944: sound1 <=  151733;
	6945: sound1 <=  173309;
	6946: sound1 <=  179108;
	6947: sound1 <=  149078;
	6948: sound1 <=  123749;
	6949: sound1 <=  105011;
	6950: sound1 <=  90393;
	6951: sound1 <=  64819;
	6952: sound1 <=  70313;
	6953: sound1 <=  54504;
	6954: sound1 <=  5920;
	6955: sound1 <=  -31830;
	6956: sound1 <=  -10681;
	6957: sound1 <=  -8881;
	6958: sound1 <=  -15503;
	6959: sound1 <=  -12878;
	6960: sound1 <=  -18524;
	6961: sound1 <=  -42236;
	6962: sound1 <=  -57281;
	6963: sound1 <=  -70374;
	6964: sound1 <=  -75470;
	6965: sound1 <=  -77789;
	6966: sound1 <=  -97015;
	6967: sound1 <=  -143585;
	6968: sound1 <=  -160950;
	6969: sound1 <=  -154999;
	6970: sound1 <=  -163513;
	6971: sound1 <=  -137848;
	6972: sound1 <=  -112854;
	6973: sound1 <=  -128021;
	6974: sound1 <=  -153198;
	6975: sound1 <=  -153809;
	6976: sound1 <=  -156555;
	6977: sound1 <=  -181946;
	6978: sound1 <=  -195343;
	6979: sound1 <=  -210388;
	6980: sound1 <=  -180725;
	6981: sound1 <=  -154968;
	6982: sound1 <=  -152954;
	6983: sound1 <=  -148254;
	6984: sound1 <=  -106415;
	6985: sound1 <=  -66254;
	6986: sound1 <=  -85297;
	6987: sound1 <=  -109955;
	6988: sound1 <=  -101501;
	6989: sound1 <=  -88806;
	6990: sound1 <=  -86792;
	6991: sound1 <=  -66040;
	6992: sound1 <=  -75043;
	6993: sound1 <=  -81238;
	6994: sound1 <=  -68390;
	6995: sound1 <=  -43640;
	6996: sound1 <=  -29755;
	6997: sound1 <=  -38666;
	6998: sound1 <=  -48676;
	6999: sound1 <=  -112091;
	7000: sound1 <=  -139526;
	7001: sound1 <=  -140961;
	7002: sound1 <=  -130035;
	7003: sound1 <=  -110168;
	7004: sound1 <=  -75745;
	7005: sound1 <=  -80505;
	7006: sound1 <=  -89203;
	7007: sound1 <=  -84503;
	7008: sound1 <=  -96191;
	7009: sound1 <=  -118713;
	7010: sound1 <=  -123993;
	7011: sound1 <=  -166443;
	7012: sound1 <=  -192474;
	7013: sound1 <=  -159943;
	7014: sound1 <=  -123413;
	7015: sound1 <=  -85480;
	7016: sound1 <=  -81146;
	7017: sound1 <=  -84717;
	7018: sound1 <=  -51086;
	7019: sound1 <=  -18524;
	7020: sound1 <=  25177;
	7021: sound1 <=  72632;
	7022: sound1 <=  96405;
	7023: sound1 <=  114380;
	7024: sound1 <=  150024;
	7025: sound1 <=  167847;
	7026: sound1 <=  190979;
	7027: sound1 <=  171692;
	7028: sound1 <=  43091;
	7029: sound1 <=  26672;
	7030: sound1 <=  7996;
	7031: sound1 <=  -37292;
	7032: sound1 <=  -43884;
	7033: sound1 <=  -51849;
	7034: sound1 <=  -59509;
	7035: sound1 <=  -30212;
	7036: sound1 <=  -9155;
	7037: sound1 <=  49652;
	7038: sound1 <=  119263;
	7039: sound1 <=  150818;
	7040: sound1 <=  176605;
	7041: sound1 <=  202850;
	7042: sound1 <=  223419;
	7043: sound1 <=  250366;
	7044: sound1 <=  289612;
	7045: sound1 <=  329590;
	7046: sound1 <=  335938;
	7047: sound1 <=  350433;
	7048: sound1 <=  354156;
	7049: sound1 <=  352478;
	7050: sound1 <=  395752;
	7051: sound1 <=  446045;
	7052: sound1 <=  389130;
	7053: sound1 <=  335541;
	7054: sound1 <=  347321;
	7055: sound1 <=  343262;
	7056: sound1 <=  361938;
	7057: sound1 <=  358154;
	7058: sound1 <=  350800;
	7059: sound1 <=  340027;
	7060: sound1 <=  333130;
	7061: sound1 <=  286957;
	7062: sound1 <=  143890;
	7063: sound1 <=  86029;
	7064: sound1 <=  74249;
	7065: sound1 <=  71259;
	7066: sound1 <=  37842;
	7067: sound1 <=  11810;
	7068: sound1 <=  20874;
	7069: sound1 <=  38391;
	7070: sound1 <=  45319;
	7071: sound1 <=  58563;
	7072: sound1 <=  91492;
	7073: sound1 <=  117981;
	7074: sound1 <=  115143;
	7075: sound1 <=  152710;
	7076: sound1 <=  200409;
	7077: sound1 <=  242218;
	7078: sound1 <=  261658;
	7079: sound1 <=  296356;
	7080: sound1 <=  235474;
	7081: sound1 <=  224091;
	7082: sound1 <=  233856;
	7083: sound1 <=  226013;
	7084: sound1 <=  236511;
	7085: sound1 <=  161163;
	7086: sound1 <=  94238;
	7087: sound1 <=  130280;
	7088: sound1 <=  122040;
	7089: sound1 <=  84320;
	7090: sound1 <=  53406;
	7091: sound1 <=  5981;
	7092: sound1 <=  -29327;
	7093: sound1 <=  -37842;
	7094: sound1 <=  -31738;
	7095: sound1 <=  -83069;
	7096: sound1 <=  -124542;
	7097: sound1 <=  -178955;
	7098: sound1 <=  -154083;
	7099: sound1 <=  -194122;
	7100: sound1 <=  -271973;
	7101: sound1 <=  -262299;
	7102: sound1 <=  -255524;
	7103: sound1 <=  -229492;
	7104: sound1 <=  -213684;
	7105: sound1 <=  -179291;
	7106: sound1 <=  -148102;
	7107: sound1 <=  -115387;
	7108: sound1 <=  -94513;
	7109: sound1 <=  -87250;
	7110: sound1 <=  -81879;
	7111: sound1 <=  -90271;
	7112: sound1 <=  -71228;
	7113: sound1 <=  -123199;
	7114: sound1 <=  -135315;
	7115: sound1 <=  -146606;
	7116: sound1 <=  -149445;
	7117: sound1 <=  -122375;
	7118: sound1 <=  -100281;
	7119: sound1 <=  -96893;
	7120: sound1 <=  -78400;
	7121: sound1 <=  -72449;
	7122: sound1 <=  -41931;
	7123: sound1 <=  -11292;
	7124: sound1 <=  14740;
	7125: sound1 <=  31952;
	7126: sound1 <=  33356;
	7127: sound1 <=  31769;
	7128: sound1 <=  42328;
	7129: sound1 <=  71350;
	7130: sound1 <=  87036;
	7131: sound1 <=  102539;
	7132: sound1 <=  109650;
	7133: sound1 <=  115448;
	7134: sound1 <=  124512;
	7135: sound1 <=  125092;
	7136: sound1 <=  127716;
	7137: sound1 <=  140106;
	7138: sound1 <=  169678;
	7139: sound1 <=  175629;
	7140: sound1 <=  174622;
	7141: sound1 <=  190460;
	7142: sound1 <=  193909;
	7143: sound1 <=  196594;
	7144: sound1 <=  160614;
	7145: sound1 <=  134827;
	7146: sound1 <=  -13275;
	7147: sound1 <=  -140747;
	7148: sound1 <=  -157135;
	7149: sound1 <=  -162628;
	7150: sound1 <=  -176453;
	7151: sound1 <=  -169617;
	7152: sound1 <=  -170319;
	7153: sound1 <=  -169464;
	7154: sound1 <=  -130219;
	7155: sound1 <=  -88104;
	7156: sound1 <=  -44098;
	7157: sound1 <=  -7172;
	7158: sound1 <=  3510;
	7159: sound1 <=  43793;
	7160: sound1 <=  88257;
	7161: sound1 <=  107697;
	7162: sound1 <=  124268;
	7163: sound1 <=  139130;
	7164: sound1 <=  160004;
	7165: sound1 <=  206665;
	7166: sound1 <=  218506;
	7167: sound1 <=  217834;
	7168: sound1 <=  243958;
	7169: sound1 <=  278931;
	7170: sound1 <=  297913;
	7171: sound1 <=  309296;
	7172: sound1 <=  310181;
	7173: sound1 <=  306976;
	7174: sound1 <=  285034;
	7175: sound1 <=  269531;
	7176: sound1 <=  259186;
	7177: sound1 <=  236267;
	7178: sound1 <=  202179;
	7179: sound1 <=  160492;
	7180: sound1 <=  124390;
	7181: sound1 <=  87402;
	7182: sound1 <=  59174;
	7183: sound1 <=  36316;
	7184: sound1 <=  -10071;
	7185: sound1 <=  -31097;
	7186: sound1 <=  -34821;
	7187: sound1 <=  -31799;
	7188: sound1 <=  -44525;
	7189: sound1 <=  -43243;
	7190: sound1 <=  -17334;
	7191: sound1 <=  -9094;
	7192: sound1 <=  -8453;
	7193: sound1 <=  11658;
	7194: sound1 <=  35217;
	7195: sound1 <=  61554;
	7196: sound1 <=  42389;
	7197: sound1 <=  35950;
	7198: sound1 <=  49896;
	7199: sound1 <=  36835;
	7200: sound1 <=  33417;
	7201: sound1 <=  28290;
	7202: sound1 <=  18372;
	7203: sound1 <=  11902;
	7204: sound1 <=  25421;
	7205: sound1 <=  4120;
	7206: sound1 <=  -40741;
	7207: sound1 <=  -43884;
	7208: sound1 <=  -39703;
	7209: sound1 <=  -61462;
	7210: sound1 <=  -65247;
	7211: sound1 <=  -81726;
	7212: sound1 <=  -122101;
	7213: sound1 <=  -142334;
	7214: sound1 <=  -186768;
	7215: sound1 <=  -210754;
	7216: sound1 <=  -195221;
	7217: sound1 <=  -193726;
	7218: sound1 <=  -187286;
	7219: sound1 <=  -161835;
	7220: sound1 <=  -160522;
	7221: sound1 <=  -167084;
	7222: sound1 <=  -150879;
	7223: sound1 <=  -134796;
	7224: sound1 <=  -125793;
	7225: sound1 <=  -103729;
	7226: sound1 <=  -91461;
	7227: sound1 <=  -125641;
	7228: sound1 <=  -180603;
	7229: sound1 <=  -213501;
	7230: sound1 <=  -252197;
	7231: sound1 <=  -283844;
	7232: sound1 <=  -273163;
	7233: sound1 <=  -254700;
	7234: sound1 <=  -255981;
	7235: sound1 <=  -251312;
	7236: sound1 <=  -256561;
	7237: sound1 <=  -238159;
	7238: sound1 <=  -229218;
	7239: sound1 <=  -239441;
	7240: sound1 <=  -220947;
	7241: sound1 <=  -194153;
	7242: sound1 <=  -187775;
	7243: sound1 <=  -177734;
	7244: sound1 <=  -165314;
	7245: sound1 <=  -159180;
	7246: sound1 <=  -158295;
	7247: sound1 <=  -144928;
	7248: sound1 <=  -127136;
	7249: sound1 <=  -101807;
	7250: sound1 <=  -60699;
	7251: sound1 <=  14130;
	7252: sound1 <=  94269;
	7253: sound1 <=  156830;
	7254: sound1 <=  204956;
	7255: sound1 <=  248199;
	7256: sound1 <=  265564;
	7257: sound1 <=  269470;
	7258: sound1 <=  252289;
	7259: sound1 <=  237946;
	7260: sound1 <=  235321;
	7261: sound1 <=  242310;
	7262: sound1 <=  212280;
	7263: sound1 <=  169098;
	7264: sound1 <=  142029;
	7265: sound1 <=  120972;
	7266: sound1 <=  127075;
	7267: sound1 <=  135040;
	7268: sound1 <=  115692;
	7269: sound1 <=  77179;
	7270: sound1 <=  51208;
	7271: sound1 <=  60516;
	7272: sound1 <=  66071;
	7273: sound1 <=  72205;
	7274: sound1 <=  81543;
	7275: sound1 <=  81879;
	7276: sound1 <=  83923;
	7277: sound1 <=  86121;
	7278: sound1 <=  103882;
	7279: sound1 <=  133942;
	7280: sound1 <=  142365;
	7281: sound1 <=  134735;
	7282: sound1 <=  158813;
	7283: sound1 <=  172852;
	7284: sound1 <=  185211;
	7285: sound1 <=  205688;
	7286: sound1 <=  222778;
	7287: sound1 <=  223175;
	7288: sound1 <=  227905;
	7289: sound1 <=  215942;
	7290: sound1 <=  188995;
	7291: sound1 <=  145386;
	7292: sound1 <=  113556;
	7293: sound1 <=  105194;
	7294: sound1 <=  83649;
	7295: sound1 <=  59692;
	7296: sound1 <=  57007;
	7297: sound1 <=  37109;
	7298: sound1 <=  6500;
	7299: sound1 <=  -3113;
	7300: sound1 <=  -20111;
	7301: sound1 <=  -132111;
	7302: sound1 <=  -156738;
	7303: sound1 <=  -185486;
	7304: sound1 <=  -188812;
	7305: sound1 <=  -136597;
	7306: sound1 <=  -100586;
	7307: sound1 <=  -89081;
	7308: sound1 <=  -62408;
	7309: sound1 <=  -17395;
	7310: sound1 <=  36163;
	7311: sound1 <=  -23712;
	7312: sound1 <=  -35004;
	7313: sound1 <=  -3052;
	7314: sound1 <=  15839;
	7315: sound1 <=  37811;
	7316: sound1 <=  37079;
	7317: sound1 <=  51270;
	7318: sound1 <=  32928;
	7319: sound1 <=  10223;
	7320: sound1 <=  -2075;
	7321: sound1 <=  -10864;
	7322: sound1 <=  -122;
	7323: sound1 <=  27527;
	7324: sound1 <=  85693;
	7325: sound1 <=  141327;
	7326: sound1 <=  68329;
	7327: sound1 <=  19257;
	7328: sound1 <=  19135;
	7329: sound1 <=  16174;
	7330: sound1 <=  29053;
	7331: sound1 <=  42633;
	7332: sound1 <=  59601;
	7333: sound1 <=  73761;
	7334: sound1 <=  75378;
	7335: sound1 <=  64331;
	7336: sound1 <=  65796;
	7337: sound1 <=  94238;
	7338: sound1 <=  121674;
	7339: sound1 <=  154633;
	7340: sound1 <=  171753;
	7341: sound1 <=  107727;
	7342: sound1 <=  129852;
	7343: sound1 <=  159058;
	7344: sound1 <=  165955;
	7345: sound1 <=  184204;
	7346: sound1 <=  171295;
	7347: sound1 <=  184692;
	7348: sound1 <=  180908;
	7349: sound1 <=  170990;
	7350: sound1 <=  156097;
	7351: sound1 <=  104736;
	7352: sound1 <=  102020;
	7353: sound1 <=  122314;
	7354: sound1 <=  122314;
	7355: sound1 <=  148529;
	7356: sound1 <=  155548;
	7357: sound1 <=  158081;
	7358: sound1 <=  188416;
	7359: sound1 <=  187683;
	7360: sound1 <=  178284;
	7361: sound1 <=  69489;
	7362: sound1 <=  8026;
	7363: sound1 <=  47333;
	7364: sound1 <=  28839;
	7365: sound1 <=  39124;
	7366: sound1 <=  32440;
	7367: sound1 <=  34058;
	7368: sound1 <=  19714;
	7369: sound1 <=  7202;
	7370: sound1 <=  23071;
	7371: sound1 <=  28595;
	7372: sound1 <=  45135;
	7373: sound1 <=  74066;
	7374: sound1 <=  34607;
	7375: sound1 <=  26978;
	7376: sound1 <=  92590;
	7377: sound1 <=  149994;
	7378: sound1 <=  191711;
	7379: sound1 <=  197601;
	7380: sound1 <=  192657;
	7381: sound1 <=  92865;
	7382: sound1 <=  68787;
	7383: sound1 <=  56854;
	7384: sound1 <=  35889;
	7385: sound1 <=  6775;
	7386: sound1 <=  -22461;
	7387: sound1 <=  -58502;
	7388: sound1 <=  -87708;
	7389: sound1 <=  -78033;
	7390: sound1 <=  -51056;
	7391: sound1 <=  -40863;
	7392: sound1 <=  -18951;
	7393: sound1 <=  12756;
	7394: sound1 <=  28961;
	7395: sound1 <=  70221;
	7396: sound1 <=  93323;
	7397: sound1 <=  136017;
	7398: sound1 <=  68237;
	7399: sound1 <=  -20752;
	7400: sound1 <=  -33478;
	7401: sound1 <=  -43671;
	7402: sound1 <=  -34790;
	7403: sound1 <=  -28015;
	7404: sound1 <=  -23682;
	7405: sound1 <=  -36896;
	7406: sound1 <=  -42114;
	7407: sound1 <=  -6897;
	7408: sound1 <=  41504;
	7409: sound1 <=  107452;
	7410: sound1 <=  150208;
	7411: sound1 <=  199799;
	7412: sound1 <=  246765;
	7413: sound1 <=  228607;
	7414: sound1 <=  209076;
	7415: sound1 <=  219757;
	7416: sound1 <=  221039;
	7417: sound1 <=  217346;
	7418: sound1 <=  178345;
	7419: sound1 <=  110077;
	7420: sound1 <=  149078;
	7421: sound1 <=  106934;
	7422: sound1 <=  90698;
	7423: sound1 <=  94696;
	7424: sound1 <=  68329;
	7425: sound1 <=  81146;
	7426: sound1 <=  74890;
	7427: sound1 <=  71533;
	7428: sound1 <=  35553;
	7429: sound1 <=  -2563;
	7430: sound1 <=  -45990;
	7431: sound1 <=  -55878;
	7432: sound1 <=  -71686;
	7433: sound1 <=  -56396;
	7434: sound1 <=  -124298;
	7435: sound1 <=  -105713;
	7436: sound1 <=  -127472;
	7437: sound1 <=  -169556;
	7438: sound1 <=  -126129;
	7439: sound1 <=  -199890;
	7440: sound1 <=  -190094;
	7441: sound1 <=  -168610;
	7442: sound1 <=  -157867;
	7443: sound1 <=  -120636;
	7444: sound1 <=  -160522;
	7445: sound1 <=  -224915;
	7446: sound1 <=  -227142;
	7447: sound1 <=  -225311;
	7448: sound1 <=  -203827;
	7449: sound1 <=  -169067;
	7450: sound1 <=  -135956;
	7451: sound1 <=  -128967;
	7452: sound1 <=  -110229;
	7453: sound1 <=  -81909;
	7454: sound1 <=  -44708;
	7455: sound1 <=  5646;
	7456: sound1 <=  60425;
	7457: sound1 <=  98694;
	7458: sound1 <=  106171;
	7459: sound1 <=  123566;
	7460: sound1 <=  153442;
	7461: sound1 <=  121002;
	7462: sound1 <=  106842;
	7463: sound1 <=  106964;
	7464: sound1 <=  108490;
	7465: sound1 <=  124512;
	7466: sound1 <=  130157;
	7467: sound1 <=  118835;
	7468: sound1 <=  99335;
	7469: sound1 <=  57465;
	7470: sound1 <=  19501;
	7471: sound1 <=  8057;
	7472: sound1 <=  -3906;
	7473: sound1 <=  16968;
	7474: sound1 <=  -132080;
	7475: sound1 <=  -249207;
	7476: sound1 <=  -265045;
	7477: sound1 <=  -293365;
	7478: sound1 <=  -307678;
	7479: sound1 <=  -307892;
	7480: sound1 <=  -278778;
	7481: sound1 <=  -233673;
	7482: sound1 <=  -199249;
	7483: sound1 <=  -160645;
	7484: sound1 <=  -120667;
	7485: sound1 <=  -52612;
	7486: sound1 <=  25787;
	7487: sound1 <=  38300;
	7488: sound1 <=  67413;
	7489: sound1 <=  97137;
	7490: sound1 <=  145050;
	7491: sound1 <=  198853;
	7492: sound1 <=  223297;
	7493: sound1 <=  234741;
	7494: sound1 <=  235565;
	7495: sound1 <=  255157;
	7496: sound1 <=  271332;
	7497: sound1 <=  288910;
	7498: sound1 <=  301056;
	7499: sound1 <=  314240;
	7500: sound1 <=  337952;
	7501: sound1 <=  339264;
	7502: sound1 <=  316803;
	7503: sound1 <=  273163;
	7504: sound1 <=  255981;
	7505: sound1 <=  248871;
	7506: sound1 <=  219574;
	7507: sound1 <=  227081;
	7508: sound1 <=  238586;
	7509: sound1 <=  216980;
	7510: sound1 <=  195190;
	7511: sound1 <=  181335;
	7512: sound1 <=  149689;
	7513: sound1 <=  136963;
	7514: sound1 <=  116364;
	7515: sound1 <=  83069;
	7516: sound1 <=  55878;
	7517: sound1 <=  45197;
	7518: sound1 <=  14435;
	7519: sound1 <=  -12573;
	7520: sound1 <=  -10406;
	7521: sound1 <=  -25269;
	7522: sound1 <=  -38666;
	7523: sound1 <=  -35980;
	7524: sound1 <=  -77728;
	7525: sound1 <=  -109650;
	7526: sound1 <=  -116638;
	7527: sound1 <=  -128784;
	7528: sound1 <=  -129425;
	7529: sound1 <=  -135529;
	7530: sound1 <=  -111359;
	7531: sound1 <=  -81543;
	7532: sound1 <=  -50964;
	7533: sound1 <=  -42603;
	7534: sound1 <=  -44647;
	7535: sound1 <=  -51880;
	7536: sound1 <=  -74310;
	7537: sound1 <=  -83710;
	7538: sound1 <=  -70587;
	7539: sound1 <=  -56854;
	7540: sound1 <=  -65521;
	7541: sound1 <=  -69214;
	7542: sound1 <=  -77545;
	7543: sound1 <=  -78186;
	7544: sound1 <=  -100281;
	7545: sound1 <=  -88593;
	7546: sound1 <=  -61737;
	7547: sound1 <=  -57892;
	7548: sound1 <=  -72632;
	7549: sound1 <=  -63507;
	7550: sound1 <=  -62103;
	7551: sound1 <=  -59875;
	7552: sound1 <=  -67535;
	7553: sound1 <=  -83954;
	7554: sound1 <=  -99762;
	7555: sound1 <=  -139923;
	7556: sound1 <=  -188751;
	7557: sound1 <=  -207092;
	7558: sound1 <=  -223114;
	7559: sound1 <=  -232208;
	7560: sound1 <=  -253113;
	7561: sound1 <=  -258911;
	7562: sound1 <=  -257294;
	7563: sound1 <=  -231720;
	7564: sound1 <=  -218658;
	7565: sound1 <=  -216125;
	7566: sound1 <=  -195038;
	7567: sound1 <=  -188721;
	7568: sound1 <=  -195465;
	7569: sound1 <=  -203674;
	7570: sound1 <=  -193542;
	7571: sound1 <=  -179810;
	7572: sound1 <=  -182159;
	7573: sound1 <=  -180145;
	7574: sound1 <=  -144135;
	7575: sound1 <=  -112091;
	7576: sound1 <=  -101379;
	7577: sound1 <=  -92682;
	7578: sound1 <=  -70190;
	7579: sound1 <=  -66162;
	7580: sound1 <=  -25024;
	7581: sound1 <=  29327;
	7582: sound1 <=  54840;
	7583: sound1 <=  114471;
	7584: sound1 <=  78339;
	7585: sound1 <=  11444;
	7586: sound1 <=  36774;
	7587: sound1 <=  47913;
	7588: sound1 <=  74127;
	7589: sound1 <=  88013;
	7590: sound1 <=  137360;
	7591: sound1 <=  139954;
	7592: sound1 <=  141205;
	7593: sound1 <=  187195;
	7594: sound1 <=  135864;
	7595: sound1 <=  171143;
	7596: sound1 <=  204102;
	7597: sound1 <=  226685;
	7598: sound1 <=  203033;
	7599: sound1 <=  229767;
	7600: sound1 <=  265778;
	7601: sound1 <=  262207;
	7602: sound1 <=  277863;
	7603: sound1 <=  295715;
	7604: sound1 <=  299866;
	7605: sound1 <=  276367;
	7606: sound1 <=  249207;
	7607: sound1 <=  226318;
	7608: sound1 <=  161438;
	7609: sound1 <=  159821;
	7610: sound1 <=  150391;
	7611: sound1 <=  175781;
	7612: sound1 <=  153503;
	7613: sound1 <=  187683;
	7614: sound1 <=  182281;
	7615: sound1 <=  131866;
	7616: sound1 <=  166199;
	7617: sound1 <=  95978;
	7618: sound1 <=  58319;
	7619: sound1 <=  104248;
	7620: sound1 <=  118774;
	7621: sound1 <=  136414;
	7622: sound1 <=  74188;
	7623: sound1 <=  82245;
	7624: sound1 <=  127014;
	7625: sound1 <=  137085;
	7626: sound1 <=  131775;
	7627: sound1 <=  128540;
	7628: sound1 <=  146027;
	7629: sound1 <=  163147;
	7630: sound1 <=  169373;
	7631: sound1 <=  197235;
	7632: sound1 <=  205933;
	7633: sound1 <=  191956;
	7634: sound1 <=  190948;
	7635: sound1 <=  193878;
	7636: sound1 <=  164337;
	7637: sound1 <=  180786;
	7638: sound1 <=  196014;
	7639: sound1 <=  178864;
	7640: sound1 <=  165741;
	7641: sound1 <=  131378;
	7642: sound1 <=  73029;
	7643: sound1 <=  142975;
	7644: sound1 <=  187073;
	7645: sound1 <=  195038;
	7646: sound1 <=  143219;
	7647: sound1 <=  87769;
	7648: sound1 <=  107391;
	7649: sound1 <=  165314;
	7650: sound1 <=  164276;
	7651: sound1 <=  82489;
	7652: sound1 <=  125793;
	7653: sound1 <=  160675;
	7654: sound1 <=  193481;
	7655: sound1 <=  177765;
	7656: sound1 <=  145172;
	7657: sound1 <=  149689;
	7658: sound1 <=  126282;
	7659: sound1 <=  36255;
	7660: sound1 <=  -27191;
	7661: sound1 <=  -6836;
	7662: sound1 <=  -1465;
	7663: sound1 <=  -74829;
	7664: sound1 <=  -66772;
	7665: sound1 <=  -116028;
	7666: sound1 <=  -149628;
	7667: sound1 <=  -97168;
	7668: sound1 <=  -85449;
	7669: sound1 <=  -24963;
	7670: sound1 <=  -22705;
	7671: sound1 <=  -35645;
	7672: sound1 <=  23743;
	7673: sound1 <=  39673;
	7674: sound1 <=  65735;
	7675: sound1 <=  76752;
	7676: sound1 <=  78522;
	7677: sound1 <=  61737;
	7678: sound1 <=  37933;
	7679: sound1 <=  -19562;
	7680: sound1 <=  -132843;
	7681: sound1 <=  -172150;
	7682: sound1 <=  -185760;
	7683: sound1 <=  -175323;
	7684: sound1 <=  -173889;
	7685: sound1 <=  -172607;
	7686: sound1 <=  -170746;
	7687: sound1 <=  -167755;
	7688: sound1 <=  -156738;
	7689: sound1 <=  -145935;
	7690: sound1 <=  -137482;
	7691: sound1 <=  -105988;
	7692: sound1 <=  -41199;
	7693: sound1 <=  1099;
	7694: sound1 <=  25665;
	7695: sound1 <=  68451;
	7696: sound1 <=  104614;
	7697: sound1 <=  131470;
	7698: sound1 <=  180389;
	7699: sound1 <=  207916;
	7700: sound1 <=  213531;
	7701: sound1 <=  236084;
	7702: sound1 <=  267578;
	7703: sound1 <=  213989;
	7704: sound1 <=  116882;
	7705: sound1 <=  123962;
	7706: sound1 <=  114380;
	7707: sound1 <=  123962;
	7708: sound1 <=  115143;
	7709: sound1 <=  88593;
	7710: sound1 <=  78735;
	7711: sound1 <=  85236;
	7712: sound1 <=  73029;
	7713: sound1 <=  53772;
	7714: sound1 <=  63324;
	7715: sound1 <=  76385;
	7716: sound1 <=  93292;
	7717: sound1 <=  126465;
	7718: sound1 <=  137573;
	7719: sound1 <=  166901;
	7720: sound1 <=  158569;
	7721: sound1 <=  152130;
	7722: sound1 <=  160950;
	7723: sound1 <=  155334;
	7724: sound1 <=  120575;
	7725: sound1 <=  16632;
	7726: sound1 <=  -107147;
	7727: sound1 <=  -145569;
	7728: sound1 <=  -196167;
	7729: sound1 <=  -226410;
	7730: sound1 <=  -212372;
	7731: sound1 <=  -185211;
	7732: sound1 <=  -175507;
	7733: sound1 <=  -187408;
	7734: sound1 <=  -138458;
	7735: sound1 <=  -77881;
	7736: sound1 <=  -97137;
	7737: sound1 <=  -52917;
	7738: sound1 <=  -19653;
	7739: sound1 <=  -8667;
	7740: sound1 <=  -97870;
	7741: sound1 <=  -141296;
	7742: sound1 <=  -112061;
	7743: sound1 <=  -77118;
	7744: sound1 <=  -79254;
	7745: sound1 <=  -77606;
	7746: sound1 <=  -83038;
	7747: sound1 <=  -85693;
	7748: sound1 <=  -78339;
	7749: sound1 <=  -61432;
	7750: sound1 <=  -71228;
	7751: sound1 <=  -96161;
	7752: sound1 <=  -122894;
	7753: sound1 <=  -127594;
	7754: sound1 <=  -98907;
	7755: sound1 <=  -50659;
	7756: sound1 <=  -41718;
	7757: sound1 <=  -61096;
	7758: sound1 <=  -35187;
	7759: sound1 <=  -21149;
	7760: sound1 <=  -27374;
	7761: sound1 <=  -42419;
	7762: sound1 <=  -66132;
	7763: sound1 <=  -77789;
	7764: sound1 <=  -77911;
	7765: sound1 <=  -83191;
	7766: sound1 <=  -91766;
	7767: sound1 <=  -109528;
	7768: sound1 <=  -121674;
	7769: sound1 <=  -116547;
	7770: sound1 <=  -101410;
	7771: sound1 <=  -169769;
	7772: sound1 <=  -220337;
	7773: sound1 <=  -212097;
	7774: sound1 <=  -202820;
	7775: sound1 <=  -187958;
	7776: sound1 <=  -167816;
	7777: sound1 <=  -120880;
	7778: sound1 <=  -114777;
	7779: sound1 <=  -102966;
	7780: sound1 <=  -49347;
	7781: sound1 <=  7751;
	7782: sound1 <=  71716;
	7783: sound1 <=  138275;
	7784: sound1 <=  204498;
	7785: sound1 <=  243713;
	7786: sound1 <=  268219;
	7787: sound1 <=  315857;
	7788: sound1 <=  370544;
	7789: sound1 <=  380127;
	7790: sound1 <=  385803;
	7791: sound1 <=  416809;
	7792: sound1 <=  446014;
	7793: sound1 <=  425079;
	7794: sound1 <=  413544;
	7795: sound1 <=  415436;
	7796: sound1 <=  424591;
	7797: sound1 <=  421417;
	7798: sound1 <=  400543;
	7799: sound1 <=  383392;
	7800: sound1 <=  377167;
	7801: sound1 <=  344727;
	7802: sound1 <=  326324;
	7803: sound1 <=  306763;
	7804: sound1 <=  279510;
	7805: sound1 <=  276306;
	7806: sound1 <=  241913;
	7807: sound1 <=  184937;
	7808: sound1 <=  68329;
	7809: sound1 <=  -101471;
	7810: sound1 <=  -180328;
	7811: sound1 <=  -230835;
	7812: sound1 <=  -273499;
	7813: sound1 <=  -309204;
	7814: sound1 <=  -326691;
	7815: sound1 <=  -326202;
	7816: sound1 <=  -298798;
	7817: sound1 <=  -274841;
	7818: sound1 <=  -258759;
	7819: sound1 <=  -241608;
	7820: sound1 <=  -219269;
	7821: sound1 <=  -217010;
	7822: sound1 <=  -206055;
	7823: sound1 <=  -161072;
	7824: sound1 <=  -146362;
	7825: sound1 <=  -146118;
	7826: sound1 <=  -139648;
	7827: sound1 <=  -117371;
	7828: sound1 <=  -100525;
	7829: sound1 <=  -78094;
	7830: sound1 <=  -48676;
	7831: sound1 <=  -26825;
	7832: sound1 <=  -27618;
	7833: sound1 <=  -23285;
	7834: sound1 <=  -6683;
	7835: sound1 <=  -28381;
	7836: sound1 <=  -31769;
	7837: sound1 <=  -33264;
	7838: sound1 <=  -18677;
	7839: sound1 <=  4089;
	7840: sound1 <=  17029;
	7841: sound1 <=  3601;
	7842: sound1 <=  -10345;
	7843: sound1 <=  -61676;
	7844: sound1 <=  -106964;
	7845: sound1 <=  -117157;
	7846: sound1 <=  -138306;
	7847: sound1 <=  -159058;
	7848: sound1 <=  -142914;
	7849: sound1 <=  -113373;
	7850: sound1 <=  -88348;
	7851: sound1 <=  -66406;
	7852: sound1 <=  -44617;
	7853: sound1 <=  -36407;
	7854: sound1 <=  -26093;
	7855: sound1 <=  2930;
	7856: sound1 <=  12329;
	7857: sound1 <=  8331;
	7858: sound1 <=  14191;
	7859: sound1 <=  45593;
	7860: sound1 <=  99701;
	7861: sound1 <=  151978;
	7862: sound1 <=  176666;
	7863: sound1 <=  166473;
	7864: sound1 <=  167480;
	7865: sound1 <=  161957;
	7866: sound1 <=  175507;
	7867: sound1 <=  176392;
	7868: sound1 <=  176239;
	7869: sound1 <=  150330;
	7870: sound1 <=  106262;
	7871: sound1 <=  102142;
	7872: sound1 <=  104736;
	7873: sound1 <=  87433;
	7874: sound1 <=  77972;
	7875: sound1 <=  76782;
	7876: sound1 <=  39764;
	7877: sound1 <=  29236;
	7878: sound1 <=  45288;
	7879: sound1 <=  50751;
	7880: sound1 <=  60547;
	7881: sound1 <=  74127;
	7882: sound1 <=  72174;
	7883: sound1 <=  59021;
	7884: sound1 <=  59052;
	7885: sound1 <=  82275;
	7886: sound1 <=  107056;
	7887: sound1 <=  123901;
	7888: sound1 <=  92773;
	7889: sound1 <=  -34485;
	7890: sound1 <=  -63965;
	7891: sound1 <=  -85266;
	7892: sound1 <=  -106262;
	7893: sound1 <=  -92010;
	7894: sound1 <=  -70160;
	7895: sound1 <=  -44952;
	7896: sound1 <=  -20996;
	7897: sound1 <=  10132;
	7898: sound1 <=  33081;
	7899: sound1 <=  54871;
	7900: sound1 <=  85968;
	7901: sound1 <=  113312;
	7902: sound1 <=  152252;
	7903: sound1 <=  197449;
	7904: sound1 <=  199829;
	7905: sound1 <=  207977;
	7906: sound1 <=  213135;
	7907: sound1 <=  210693;
	7908: sound1 <=  216644;
	7909: sound1 <=  224304;
	7910: sound1 <=  234467;
	7911: sound1 <=  216095;
	7912: sound1 <=  221985;
	7913: sound1 <=  254028;
	7914: sound1 <=  268341;
	7915: sound1 <=  286499;
	7916: sound1 <=  283508;
	7917: sound1 <=  262543;
	7918: sound1 <=  283173;
	7919: sound1 <=  311920;
	7920: sound1 <=  355957;
	7921: sound1 <=  358459;
	7922: sound1 <=  345612;
	7923: sound1 <=  324585;
	7924: sound1 <=  290222;
	7925: sound1 <=  257446;
	7926: sound1 <=  220520;
	7927: sound1 <=  187012;
	7928: sound1 <=  177826;
	7929: sound1 <=  171783;
	7930: sound1 <=  156647;
	7931: sound1 <=  158417;
	7932: sound1 <=  157715;
	7933: sound1 <=  158325;
	7934: sound1 <=  169952;
	7935: sound1 <=  169495;
	7936: sound1 <=  153076;
	7937: sound1 <=  124512;
	7938: sound1 <=  110779;
	7939: sound1 <=  123077;
	7940: sound1 <=  124542;
	7941: sound1 <=  81879;
	7942: sound1 <=  52155;
	7943: sound1 <=  25330;
	7944: sound1 <=  -7782;
	7945: sound1 <=  -54596;
	7946: sound1 <=  -106781;
	7947: sound1 <=  -174042;
	7948: sound1 <=  -207092;
	7949: sound1 <=  -261108;
	7950: sound1 <=  -323486;
	7951: sound1 <=  -355927;
	7952: sound1 <=  -345520;
	7953: sound1 <=  -330566;
	7954: sound1 <=  -323090;
	7955: sound1 <=  -316376;
	7956: sound1 <=  -324341;
	7957: sound1 <=  -315796;
	7958: sound1 <=  -308929;
	7959: sound1 <=  -297516;
	7960: sound1 <=  -270599;
	7961: sound1 <=  -274506;
	7962: sound1 <=  -288086;
	7963: sound1 <=  -273499;
	7964: sound1 <=  -227814;
	7965: sound1 <=  -180725;
	7966: sound1 <=  -151276;
	7967: sound1 <=  -109528;
	7968: sound1 <=  -65857;
	7969: sound1 <=  -58075;
	7970: sound1 <=  -31128;
	7971: sound1 <=  3845;
	7972: sound1 <=  28198;
	7973: sound1 <=  46783;
	7974: sound1 <=  38483;
	7975: sound1 <=  35583;
	7976: sound1 <=  42389;
	7977: sound1 <=  36530;
	7978: sound1 <=  23895;
	7979: sound1 <=  -30243;
	7980: sound1 <=  -41351;
	7981: sound1 <=  -85632;
	7982: sound1 <=  -122803;
	7983: sound1 <=  -114258;
	7984: sound1 <=  -88013;
	7985: sound1 <=  -98419;
	7986: sound1 <=  -115143;
	7987: sound1 <=  -129089;
	7988: sound1 <=  -128754;
	7989: sound1 <=  -109741;
	7990: sound1 <=  -93903;
	7991: sound1 <=  -74036;
	7992: sound1 <=  -58899;
	7993: sound1 <=  -66498;
	7994: sound1 <=  -76355;
	7995: sound1 <=  -53772;
	7996: sound1 <=  -20447;
	7997: sound1 <=  732;
	7998: sound1 <=  9674;
	7999: sound1 <=  32013;
	8000: sound1 <=  69427;
	8001: sound1 <=  124756;
	8002: sound1 <=  171326;
	8003: sound1 <=  202637;
	8004: sound1 <=  221954;
	8005: sound1 <=  208344;
	8006: sound1 <=  215881;
	8007: sound1 <=  131287;
	8008: sound1 <=  -7813;
	8009: sound1 <=  -44250;
	8010: sound1 <=  -76721;
	8011: sound1 <=  -80292;
	8012: sound1 <=  -62744;
	8013: sound1 <=  -36804;
	8014: sound1 <=  -58655;
	8015: sound1 <=  -47791;
	8016: sound1 <=  -9003;
	8017: sound1 <=  8484;
	8018: sound1 <=  15442;
	8019: sound1 <=  19318;
	8020: sound1 <=  49957;
	8021: sound1 <=  108826;
	8022: sound1 <=  154449;
	8023: sound1 <=  184235;
	8024: sound1 <=  203217;
	8025: sound1 <=  211884;
	8026: sound1 <=  241669;
	8027: sound1 <=  261108;
	8028: sound1 <=  268311;
	8029: sound1 <=  285950;
	8030: sound1 <=  286713;
	8031: sound1 <=  285461;
	8032: sound1 <=  283691;
	8033: sound1 <=  290771;
	8034: sound1 <=  291626;
	8035: sound1 <=  297424;
	8036: sound1 <=  326904;
	8037: sound1 <=  340271;
	8038: sound1 <=  220825;
	8039: sound1 <=  131836;
	8040: sound1 <=  86853;
	8041: sound1 <=  37201;
	8042: sound1 <=  -13245;
	8043: sound1 <=  -42053;
	8044: sound1 <=  -54688;
	8045: sound1 <=  -77393;
	8046: sound1 <=  -116486;
	8047: sound1 <=  -152832;
	8048: sound1 <=  -157104;
	8049: sound1 <=  -155334;
	8050: sound1 <=  -152588;
	8051: sound1 <=  -157715;
	8052: sound1 <=  -157135;
	8053: sound1 <=  -97687;
	8054: sound1 <=  -32074;
	8055: sound1 <=  366;
	8056: sound1 <=  60822;
	8057: sound1 <=  120605;
	8058: sound1 <=  154266;
	8059: sound1 <=  216339;
	8060: sound1 <=  247559;
	8061: sound1 <=  270447;
	8062: sound1 <=  291504;
	8063: sound1 <=  264343;
	8064: sound1 <=  253052;
	8065: sound1 <=  241730;
	8066: sound1 <=  234375;
	8067: sound1 <=  265259;
	8068: sound1 <=  281769;
	8069: sound1 <=  279877;
	8070: sound1 <=  253815;
	8071: sound1 <=  230194;
	8072: sound1 <=  230255;
	8073: sound1 <=  210358;
	8074: sound1 <=  169586;
	8075: sound1 <=  145233;
	8076: sound1 <=  130280;
	8077: sound1 <=  116089;
	8078: sound1 <=  101898;
	8079: sound1 <=  75531;
	8080: sound1 <=  47119;
	8081: sound1 <=  20599;
	8082: sound1 <=  -15869;
	8083: sound1 <=  -42267;
	8084: sound1 <=  -109802;
	8085: sound1 <=  -156952;
	8086: sound1 <=  -178772;
	8087: sound1 <=  -201965;
	8088: sound1 <=  -196777;
	8089: sound1 <=  -154907;
	8090: sound1 <=  -128815;
	8091: sound1 <=  -122650;
	8092: sound1 <=  -122833;
	8093: sound1 <=  -105621;
	8094: sound1 <=  -90973;
	8095: sound1 <=  -79224;
	8096: sound1 <=  -44769;
	8097: sound1 <=  -47791;
	8098: sound1 <=  -57465;
	8099: sound1 <=  -42694;
	8100: sound1 <=  -23712;
	8101: sound1 <=  5096;
	8102: sound1 <=  54199;
	8103: sound1 <=  51208;
	8104: sound1 <=  75989;
	8105: sound1 <=  100250;
	8106: sound1 <=  90485;
	8107: sound1 <=  90729;
	8108: sound1 <=  70099;
	8109: sound1 <=  51086;
	8110: sound1 <=  18158;
	8111: sound1 <=  -17975;
	8112: sound1 <=  -19897;
	8113: sound1 <=  -12238;
	8114: sound1 <=  -18555;
	8115: sound1 <=  -23438;
	8116: sound1 <=  -34760;
	8117: sound1 <=  -46173;
	8118: sound1 <=  -47241;
	8119: sound1 <=  -46051;
	8120: sound1 <=  -62408;
	8121: sound1 <=  -51697;
	8122: sound1 <=  -85419;
	8123: sound1 <=  -200897;
	8124: sound1 <=  -210693;
	8125: sound1 <=  -200714;
	8126: sound1 <=  -202423;
	8127: sound1 <=  -212402;
	8128: sound1 <=  -221252;
	8129: sound1 <=  -217743;
	8130: sound1 <=  -196777;
	8131: sound1 <=  -148621;
	8132: sound1 <=  -134827;
	8133: sound1 <=  -127167;
	8134: sound1 <=  -86060;
	8135: sound1 <=  -58258;
	8136: sound1 <=  -43304;
	8137: sound1 <=  -76477;
	8138: sound1 <=  -54413;
	8139: sound1 <=  -19012;
	8140: sound1 <=  23010;
	8141: sound1 <=  74677;
	8142: sound1 <=  50751;
	8143: sound1 <=  41595;
	8144: sound1 <=  93872;
	8145: sound1 <=  140198;
	8146: sound1 <=  108826;
	8147: sound1 <=  72571;
	8148: sound1 <=  71686;
	8149: sound1 <=  58014;
	8150: sound1 <=  63324;
	8151: sound1 <=  77271;
	8152: sound1 <=  73334;
	8153: sound1 <=  82642;
	8154: sound1 <=  92682;
	8155: sound1 <=  94269;
	8156: sound1 <=  100098;
	8157: sound1 <=  118317;
	8158: sound1 <=  132629;
	8159: sound1 <=  139923;
	8160: sound1 <=  134399;
	8161: sound1 <=  150665;
	8162: sound1 <=  149078;
	8163: sound1 <=  108368;
	8164: sound1 <=  79376;
	8165: sound1 <=  81207;
	8166: sound1 <=  99182;
	8167: sound1 <=  111237;
	8168: sound1 <=  81055;
	8169: sound1 <=  -34668;
	8170: sound1 <=  -84351;
	8171: sound1 <=  -79529;
	8172: sound1 <=  -52673;
	8173: sound1 <=  -59601;
	8174: sound1 <=  -32654;
	8175: sound1 <=  6958;
	8176: sound1 <=  17883;
	8177: sound1 <=  32074;
	8178: sound1 <=  25269;
	8179: sound1 <=  35492;
	8180: sound1 <=  70862;
	8181: sound1 <=  106720;
	8182: sound1 <=  128571;
	8183: sound1 <=  144135;
	8184: sound1 <=  164764;
	8185: sound1 <=  198730;
	8186: sound1 <=  199402;
	8187: sound1 <=  207397;
	8188: sound1 <=  222473;
	8189: sound1 <=  243378;
	8190: sound1 <=  251465;
	8191: begin
				sound1 <=  244781;
				start <= 1'b0;
				testi <= 1'b0;
			end

	default: sound1 <= 0;
endcase
		
		
		
	end else delay_cnt <= delay_cnt + 17'd1;
	end
end

/*****************************************************************************
 *                            Combinational Logic                            *
 *****************************************************************************/

//assign delay = {SW[3:0], 15'd3000};

wire [31:0] sound = (test == 0) ? 0 : 500*sound1;
wire test = testi;

assign read_audio_in			= audio_in_available & audio_out_allowed;

assign left_channel_audio_out	= left_channel_audio_in+sound;
assign right_channel_audio_out	= right_channel_audio_in+sound;
assign write_audio_out			= audio_in_available & audio_out_allowed;

/*****************************************************************************
 *                              Internal Modules                             *
 *****************************************************************************/

Audio_Controller Audio_Controller (
	// Inputs
	.CLOCK_50						(CLOCK_50),
	.reset						(~KEY[0]),

	.clear_audio_in_memory		(),
	.read_audio_in				(read_audio_in),
	
	.clear_audio_out_memory		(),
	.left_channel_audio_out		(left_channel_audio_out),
	.right_channel_audio_out	(right_channel_audio_out),
	.write_audio_out			(write_audio_out),

	.AUD_ADCDAT					(AUD_ADCDAT),

	// Bidirectionals
	.AUD_BCLK					(AUD_BCLK),
	.AUD_ADCLRCK				(AUD_ADCLRCK),
	.AUD_DACLRCK				(AUD_DACLRCK),


	// Outputs
	.audio_in_available			(audio_in_available),
	.left_channel_audio_in		(left_channel_audio_in),
	.right_channel_audio_in		(right_channel_audio_in),

	.audio_out_allowed			(audio_out_allowed),

	.AUD_XCK					(AUD_XCK),
	.AUD_DACDAT					(AUD_DACDAT)

);

avconf #(.USE_MIC_INPUT(1)) avc (
	.I2C_SCLK					(I2C_SCLK),
	.I2C_SDAT					(I2C_SDAT),
	.CLOCK_50					(CLOCK_50),
	.reset						(~KEY[0])
);

endmodule

